`ifndef __COMMON_OFDM_VH__
	`define __COMMON_OFDM_VH__

//parameter	DATA_FFT_SIZE = 16;
//parameter	DATA_FFT_FAST_SIZE = 16;

`define PILOT_P13_I      1024
`define PILOT_P38_I      1024
`define PILOT_P63_I      1024
`define PILOT_P88_I      1024
`define PILOT_P_88_I     1024
`define PILOT_P_63_I     1024
`define PILOT_P_38_I     1024
`define PILOT_P_13_I     1024

`define PILOT_P13_Q      1024
`define PILOT_P38_Q      1024
`define PILOT_P63_Q      1024
`define PILOT_P88_Q      1024
`define PILOT_P_88_Q     1024
`define PILOT_P_63_Q     1024
`define PILOT_P_38_Q     1024
`define PILOT_P_13_Q     1024

`endif //__COMMON_OFDM_VH__