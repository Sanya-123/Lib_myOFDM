`ifndef __COMMON_VH__
	`define __COMMON_VH__

parameter	DATA_FFT_SIZE = 16;
parameter	DATA_FFT_FAST_SIZE = 16;

`endif //__COMMON_VH__