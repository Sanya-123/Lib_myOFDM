module dds_romb
  (
  iclk    ,
  iclkena ,
  iadr0   ,
  iadr1   ,
  odat0   ,
  odat1
  );

  input               iclk;
  input               iclkena;
  input        [12:0] iadr0;
  input        [12:0] iadr1;
  output logic [12:0] odat0;
  output logic [12:0] odat1;

  localparam bit [12:0] coe [0:8191] = '{
      0 ,    // 0
      2 ,    // 1
      3 ,    // 2
      5 ,    // 3
      6 ,    // 4
      8 ,    // 5
      9 ,    // 6
      11 ,    // 7
      13 ,    // 8
      14 ,    // 9
      16 ,    // 10
      17 ,    // 11
      19 ,    // 12
      20 ,    // 13
      22 ,    // 14
      24 ,    // 15
      25 ,    // 16
      27 ,    // 17
      28 ,    // 18
      30 ,    // 19
      31 ,    // 20
      33 ,    // 21
      35 ,    // 22
      36 ,    // 23
      38 ,    // 24
      39 ,    // 25
      41 ,    // 26
      42 ,    // 27
      44 ,    // 28
      45 ,    // 29
      47 ,    // 30
      49 ,    // 31
      50 ,    // 32
      52 ,    // 33
      53 ,    // 34
      55 ,    // 35
      56 ,    // 36
      58 ,    // 37
      60 ,    // 38
      61 ,    // 39
      63 ,    // 40
      64 ,    // 41
      66 ,    // 42
      67 ,    // 43
      69 ,    // 44
      71 ,    // 45
      72 ,    // 46
      74 ,    // 47
      75 ,    // 48
      77 ,    // 49
      78 ,    // 50
      80 ,    // 51
      82 ,    // 52
      83 ,    // 53
      85 ,    // 54
      86 ,    // 55
      88 ,    // 56
      89 ,    // 57
      91 ,    // 58
      93 ,    // 59
      94 ,    // 60
      96 ,    // 61
      97 ,    // 62
      99 ,    // 63
      100 ,    // 64
      102 ,    // 65
      104 ,    // 66
      105 ,    // 67
      107 ,    // 68
      108 ,    // 69
      110 ,    // 70
      111 ,    // 71
      113 ,    // 72
      115 ,    // 73
      116 ,    // 74
      118 ,    // 75
      119 ,    // 76
      121 ,    // 77
      122 ,    // 78
      124 ,    // 79
      125 ,    // 80
      127 ,    // 81
      129 ,    // 82
      130 ,    // 83
      132 ,    // 84
      133 ,    // 85
      135 ,    // 86
      136 ,    // 87
      138 ,    // 88
      140 ,    // 89
      141 ,    // 90
      143 ,    // 91
      144 ,    // 92
      146 ,    // 93
      147 ,    // 94
      149 ,    // 95
      151 ,    // 96
      152 ,    // 97
      154 ,    // 98
      155 ,    // 99
      157 ,    // 100
      158 ,    // 101
      160 ,    // 102
      162 ,    // 103
      163 ,    // 104
      165 ,    // 105
      166 ,    // 106
      168 ,    // 107
      169 ,    // 108
      171 ,    // 109
      173 ,    // 110
      174 ,    // 111
      176 ,    // 112
      177 ,    // 113
      179 ,    // 114
      180 ,    // 115
      182 ,    // 116
      184 ,    // 117
      185 ,    // 118
      187 ,    // 119
      188 ,    // 120
      190 ,    // 121
      191 ,    // 122
      193 ,    // 123
      195 ,    // 124
      196 ,    // 125
      198 ,    // 126
      199 ,    // 127
      201 ,    // 128
      202 ,    // 129
      204 ,    // 130
      205 ,    // 131
      207 ,    // 132
      209 ,    // 133
      210 ,    // 134
      212 ,    // 135
      213 ,    // 136
      215 ,    // 137
      216 ,    // 138
      218 ,    // 139
      220 ,    // 140
      221 ,    // 141
      223 ,    // 142
      224 ,    // 143
      226 ,    // 144
      227 ,    // 145
      229 ,    // 146
      231 ,    // 147
      232 ,    // 148
      234 ,    // 149
      235 ,    // 150
      237 ,    // 151
      238 ,    // 152
      240 ,    // 153
      242 ,    // 154
      243 ,    // 155
      245 ,    // 156
      246 ,    // 157
      248 ,    // 158
      249 ,    // 159
      251 ,    // 160
      253 ,    // 161
      254 ,    // 162
      256 ,    // 163
      257 ,    // 164
      259 ,    // 165
      260 ,    // 166
      262 ,    // 167
      263 ,    // 168
      265 ,    // 169
      267 ,    // 170
      268 ,    // 171
      270 ,    // 172
      271 ,    // 173
      273 ,    // 174
      274 ,    // 175
      276 ,    // 176
      278 ,    // 177
      279 ,    // 178
      281 ,    // 179
      282 ,    // 180
      284 ,    // 181
      285 ,    // 182
      287 ,    // 183
      289 ,    // 184
      290 ,    // 185
      292 ,    // 186
      293 ,    // 187
      295 ,    // 188
      296 ,    // 189
      298 ,    // 190
      300 ,    // 191
      301 ,    // 192
      303 ,    // 193
      304 ,    // 194
      306 ,    // 195
      307 ,    // 196
      309 ,    // 197
      311 ,    // 198
      312 ,    // 199
      314 ,    // 200
      315 ,    // 201
      317 ,    // 202
      318 ,    // 203
      320 ,    // 204
      322 ,    // 205
      323 ,    // 206
      325 ,    // 207
      326 ,    // 208
      328 ,    // 209
      329 ,    // 210
      331 ,    // 211
      332 ,    // 212
      334 ,    // 213
      336 ,    // 214
      337 ,    // 215
      339 ,    // 216
      340 ,    // 217
      342 ,    // 218
      343 ,    // 219
      345 ,    // 220
      347 ,    // 221
      348 ,    // 222
      350 ,    // 223
      351 ,    // 224
      353 ,    // 225
      354 ,    // 226
      356 ,    // 227
      358 ,    // 228
      359 ,    // 229
      361 ,    // 230
      362 ,    // 231
      364 ,    // 232
      365 ,    // 233
      367 ,    // 234
      369 ,    // 235
      370 ,    // 236
      372 ,    // 237
      373 ,    // 238
      375 ,    // 239
      376 ,    // 240
      378 ,    // 241
      379 ,    // 242
      381 ,    // 243
      383 ,    // 244
      384 ,    // 245
      386 ,    // 246
      387 ,    // 247
      389 ,    // 248
      390 ,    // 249
      392 ,    // 250
      394 ,    // 251
      395 ,    // 252
      397 ,    // 253
      398 ,    // 254
      400 ,    // 255
      401 ,    // 256
      403 ,    // 257
      405 ,    // 258
      406 ,    // 259
      408 ,    // 260
      409 ,    // 261
      411 ,    // 262
      412 ,    // 263
      414 ,    // 264
      416 ,    // 265
      417 ,    // 266
      419 ,    // 267
      420 ,    // 268
      422 ,    // 269
      423 ,    // 270
      425 ,    // 271
      426 ,    // 272
      428 ,    // 273
      430 ,    // 274
      431 ,    // 275
      433 ,    // 276
      434 ,    // 277
      436 ,    // 278
      437 ,    // 279
      439 ,    // 280
      441 ,    // 281
      442 ,    // 282
      444 ,    // 283
      445 ,    // 284
      447 ,    // 285
      448 ,    // 286
      450 ,    // 287
      452 ,    // 288
      453 ,    // 289
      455 ,    // 290
      456 ,    // 291
      458 ,    // 292
      459 ,    // 293
      461 ,    // 294
      463 ,    // 295
      464 ,    // 296
      466 ,    // 297
      467 ,    // 298
      469 ,    // 299
      470 ,    // 300
      472 ,    // 301
      473 ,    // 302
      475 ,    // 303
      477 ,    // 304
      478 ,    // 305
      480 ,    // 306
      481 ,    // 307
      483 ,    // 308
      484 ,    // 309
      486 ,    // 310
      488 ,    // 311
      489 ,    // 312
      491 ,    // 313
      492 ,    // 314
      494 ,    // 315
      495 ,    // 316
      497 ,    // 317
      499 ,    // 318
      500 ,    // 319
      502 ,    // 320
      503 ,    // 321
      505 ,    // 322
      506 ,    // 323
      508 ,    // 324
      509 ,    // 325
      511 ,    // 326
      513 ,    // 327
      514 ,    // 328
      516 ,    // 329
      517 ,    // 330
      519 ,    // 331
      520 ,    // 332
      522 ,    // 333
      524 ,    // 334
      525 ,    // 335
      527 ,    // 336
      528 ,    // 337
      530 ,    // 338
      531 ,    // 339
      533 ,    // 340
      535 ,    // 341
      536 ,    // 342
      538 ,    // 343
      539 ,    // 344
      541 ,    // 345
      542 ,    // 346
      544 ,    // 347
      546 ,    // 348
      547 ,    // 349
      549 ,    // 350
      550 ,    // 351
      552 ,    // 352
      553 ,    // 353
      555 ,    // 354
      556 ,    // 355
      558 ,    // 356
      560 ,    // 357
      561 ,    // 358
      563 ,    // 359
      564 ,    // 360
      566 ,    // 361
      567 ,    // 362
      569 ,    // 363
      571 ,    // 364
      572 ,    // 365
      574 ,    // 366
      575 ,    // 367
      577 ,    // 368
      578 ,    // 369
      580 ,    // 370
      581 ,    // 371
      583 ,    // 372
      585 ,    // 373
      586 ,    // 374
      588 ,    // 375
      589 ,    // 376
      591 ,    // 377
      592 ,    // 378
      594 ,    // 379
      596 ,    // 380
      597 ,    // 381
      599 ,    // 382
      600 ,    // 383
      602 ,    // 384
      603 ,    // 385
      605 ,    // 386
      607 ,    // 387
      608 ,    // 388
      610 ,    // 389
      611 ,    // 390
      613 ,    // 391
      614 ,    // 392
      616 ,    // 393
      617 ,    // 394
      619 ,    // 395
      621 ,    // 396
      622 ,    // 397
      624 ,    // 398
      625 ,    // 399
      627 ,    // 400
      628 ,    // 401
      630 ,    // 402
      632 ,    // 403
      633 ,    // 404
      635 ,    // 405
      636 ,    // 406
      638 ,    // 407
      639 ,    // 408
      641 ,    // 409
      643 ,    // 410
      644 ,    // 411
      646 ,    // 412
      647 ,    // 413
      649 ,    // 414
      650 ,    // 415
      652 ,    // 416
      653 ,    // 417
      655 ,    // 418
      657 ,    // 419
      658 ,    // 420
      660 ,    // 421
      661 ,    // 422
      663 ,    // 423
      664 ,    // 424
      666 ,    // 425
      668 ,    // 426
      669 ,    // 427
      671 ,    // 428
      672 ,    // 429
      674 ,    // 430
      675 ,    // 431
      677 ,    // 432
      678 ,    // 433
      680 ,    // 434
      682 ,    // 435
      683 ,    // 436
      685 ,    // 437
      686 ,    // 438
      688 ,    // 439
      689 ,    // 440
      691 ,    // 441
      693 ,    // 442
      694 ,    // 443
      696 ,    // 444
      697 ,    // 445
      699 ,    // 446
      700 ,    // 447
      702 ,    // 448
      703 ,    // 449
      705 ,    // 450
      707 ,    // 451
      708 ,    // 452
      710 ,    // 453
      711 ,    // 454
      713 ,    // 455
      714 ,    // 456
      716 ,    // 457
      718 ,    // 458
      719 ,    // 459
      721 ,    // 460
      722 ,    // 461
      724 ,    // 462
      725 ,    // 463
      727 ,    // 464
      728 ,    // 465
      730 ,    // 466
      732 ,    // 467
      733 ,    // 468
      735 ,    // 469
      736 ,    // 470
      738 ,    // 471
      739 ,    // 472
      741 ,    // 473
      743 ,    // 474
      744 ,    // 475
      746 ,    // 476
      747 ,    // 477
      749 ,    // 478
      750 ,    // 479
      752 ,    // 480
      753 ,    // 481
      755 ,    // 482
      757 ,    // 483
      758 ,    // 484
      760 ,    // 485
      761 ,    // 486
      763 ,    // 487
      764 ,    // 488
      766 ,    // 489
      768 ,    // 490
      769 ,    // 491
      771 ,    // 492
      772 ,    // 493
      774 ,    // 494
      775 ,    // 495
      777 ,    // 496
      778 ,    // 497
      780 ,    // 498
      782 ,    // 499
      783 ,    // 500
      785 ,    // 501
      786 ,    // 502
      788 ,    // 503
      789 ,    // 504
      791 ,    // 505
      793 ,    // 506
      794 ,    // 507
      796 ,    // 508
      797 ,    // 509
      799 ,    // 510
      800 ,    // 511
      802 ,    // 512
      803 ,    // 513
      805 ,    // 514
      807 ,    // 515
      808 ,    // 516
      810 ,    // 517
      811 ,    // 518
      813 ,    // 519
      814 ,    // 520
      816 ,    // 521
      817 ,    // 522
      819 ,    // 523
      821 ,    // 524
      822 ,    // 525
      824 ,    // 526
      825 ,    // 527
      827 ,    // 528
      828 ,    // 529
      830 ,    // 530
      832 ,    // 531
      833 ,    // 532
      835 ,    // 533
      836 ,    // 534
      838 ,    // 535
      839 ,    // 536
      841 ,    // 537
      842 ,    // 538
      844 ,    // 539
      846 ,    // 540
      847 ,    // 541
      849 ,    // 542
      850 ,    // 543
      852 ,    // 544
      853 ,    // 545
      855 ,    // 546
      857 ,    // 547
      858 ,    // 548
      860 ,    // 549
      861 ,    // 550
      863 ,    // 551
      864 ,    // 552
      866 ,    // 553
      867 ,    // 554
      869 ,    // 555
      871 ,    // 556
      872 ,    // 557
      874 ,    // 558
      875 ,    // 559
      877 ,    // 560
      878 ,    // 561
      880 ,    // 562
      881 ,    // 563
      883 ,    // 564
      885 ,    // 565
      886 ,    // 566
      888 ,    // 567
      889 ,    // 568
      891 ,    // 569
      892 ,    // 570
      894 ,    // 571
      895 ,    // 572
      897 ,    // 573
      899 ,    // 574
      900 ,    // 575
      902 ,    // 576
      903 ,    // 577
      905 ,    // 578
      906 ,    // 579
      908 ,    // 580
      910 ,    // 581
      911 ,    // 582
      913 ,    // 583
      914 ,    // 584
      916 ,    // 585
      917 ,    // 586
      919 ,    // 587
      920 ,    // 588
      922 ,    // 589
      924 ,    // 590
      925 ,    // 591
      927 ,    // 592
      928 ,    // 593
      930 ,    // 594
      931 ,    // 595
      933 ,    // 596
      934 ,    // 597
      936 ,    // 598
      938 ,    // 599
      939 ,    // 600
      941 ,    // 601
      942 ,    // 602
      944 ,    // 603
      945 ,    // 604
      947 ,    // 605
      948 ,    // 606
      950 ,    // 607
      952 ,    // 608
      953 ,    // 609
      955 ,    // 610
      956 ,    // 611
      958 ,    // 612
      959 ,    // 613
      961 ,    // 614
      963 ,    // 615
      964 ,    // 616
      966 ,    // 617
      967 ,    // 618
      969 ,    // 619
      970 ,    // 620
      972 ,    // 621
      973 ,    // 622
      975 ,    // 623
      977 ,    // 624
      978 ,    // 625
      980 ,    // 626
      981 ,    // 627
      983 ,    // 628
      984 ,    // 629
      986 ,    // 630
      987 ,    // 631
      989 ,    // 632
      991 ,    // 633
      992 ,    // 634
      994 ,    // 635
      995 ,    // 636
      997 ,    // 637
      998 ,    // 638
      1000 ,    // 639
      1001 ,    // 640
      1003 ,    // 641
      1005 ,    // 642
      1006 ,    // 643
      1008 ,    // 644
      1009 ,    // 645
      1011 ,    // 646
      1012 ,    // 647
      1014 ,    // 648
      1015 ,    // 649
      1017 ,    // 650
      1019 ,    // 651
      1020 ,    // 652
      1022 ,    // 653
      1023 ,    // 654
      1025 ,    // 655
      1026 ,    // 656
      1028 ,    // 657
      1029 ,    // 658
      1031 ,    // 659
      1033 ,    // 660
      1034 ,    // 661
      1036 ,    // 662
      1037 ,    // 663
      1039 ,    // 664
      1040 ,    // 665
      1042 ,    // 666
      1043 ,    // 667
      1045 ,    // 668
      1047 ,    // 669
      1048 ,    // 670
      1050 ,    // 671
      1051 ,    // 672
      1053 ,    // 673
      1054 ,    // 674
      1056 ,    // 675
      1057 ,    // 676
      1059 ,    // 677
      1061 ,    // 678
      1062 ,    // 679
      1064 ,    // 680
      1065 ,    // 681
      1067 ,    // 682
      1068 ,    // 683
      1070 ,    // 684
      1071 ,    // 685
      1073 ,    // 686
      1075 ,    // 687
      1076 ,    // 688
      1078 ,    // 689
      1079 ,    // 690
      1081 ,    // 691
      1082 ,    // 692
      1084 ,    // 693
      1085 ,    // 694
      1087 ,    // 695
      1089 ,    // 696
      1090 ,    // 697
      1092 ,    // 698
      1093 ,    // 699
      1095 ,    // 700
      1096 ,    // 701
      1098 ,    // 702
      1099 ,    // 703
      1101 ,    // 704
      1103 ,    // 705
      1104 ,    // 706
      1106 ,    // 707
      1107 ,    // 708
      1109 ,    // 709
      1110 ,    // 710
      1112 ,    // 711
      1113 ,    // 712
      1115 ,    // 713
      1117 ,    // 714
      1118 ,    // 715
      1120 ,    // 716
      1121 ,    // 717
      1123 ,    // 718
      1124 ,    // 719
      1126 ,    // 720
      1127 ,    // 721
      1129 ,    // 722
      1131 ,    // 723
      1132 ,    // 724
      1134 ,    // 725
      1135 ,    // 726
      1137 ,    // 727
      1138 ,    // 728
      1140 ,    // 729
      1141 ,    // 730
      1143 ,    // 731
      1145 ,    // 732
      1146 ,    // 733
      1148 ,    // 734
      1149 ,    // 735
      1151 ,    // 736
      1152 ,    // 737
      1154 ,    // 738
      1155 ,    // 739
      1157 ,    // 740
      1158 ,    // 741
      1160 ,    // 742
      1162 ,    // 743
      1163 ,    // 744
      1165 ,    // 745
      1166 ,    // 746
      1168 ,    // 747
      1169 ,    // 748
      1171 ,    // 749
      1172 ,    // 750
      1174 ,    // 751
      1176 ,    // 752
      1177 ,    // 753
      1179 ,    // 754
      1180 ,    // 755
      1182 ,    // 756
      1183 ,    // 757
      1185 ,    // 758
      1186 ,    // 759
      1188 ,    // 760
      1190 ,    // 761
      1191 ,    // 762
      1193 ,    // 763
      1194 ,    // 764
      1196 ,    // 765
      1197 ,    // 766
      1199 ,    // 767
      1200 ,    // 768
      1202 ,    // 769
      1204 ,    // 770
      1205 ,    // 771
      1207 ,    // 772
      1208 ,    // 773
      1210 ,    // 774
      1211 ,    // 775
      1213 ,    // 776
      1214 ,    // 777
      1216 ,    // 778
      1217 ,    // 779
      1219 ,    // 780
      1221 ,    // 781
      1222 ,    // 782
      1224 ,    // 783
      1225 ,    // 784
      1227 ,    // 785
      1228 ,    // 786
      1230 ,    // 787
      1231 ,    // 788
      1233 ,    // 789
      1235 ,    // 790
      1236 ,    // 791
      1238 ,    // 792
      1239 ,    // 793
      1241 ,    // 794
      1242 ,    // 795
      1244 ,    // 796
      1245 ,    // 797
      1247 ,    // 798
      1248 ,    // 799
      1250 ,    // 800
      1252 ,    // 801
      1253 ,    // 802
      1255 ,    // 803
      1256 ,    // 804
      1258 ,    // 805
      1259 ,    // 806
      1261 ,    // 807
      1262 ,    // 808
      1264 ,    // 809
      1266 ,    // 810
      1267 ,    // 811
      1269 ,    // 812
      1270 ,    // 813
      1272 ,    // 814
      1273 ,    // 815
      1275 ,    // 816
      1276 ,    // 817
      1278 ,    // 818
      1279 ,    // 819
      1281 ,    // 820
      1283 ,    // 821
      1284 ,    // 822
      1286 ,    // 823
      1287 ,    // 824
      1289 ,    // 825
      1290 ,    // 826
      1292 ,    // 827
      1293 ,    // 828
      1295 ,    // 829
      1297 ,    // 830
      1298 ,    // 831
      1300 ,    // 832
      1301 ,    // 833
      1303 ,    // 834
      1304 ,    // 835
      1306 ,    // 836
      1307 ,    // 837
      1309 ,    // 838
      1310 ,    // 839
      1312 ,    // 840
      1314 ,    // 841
      1315 ,    // 842
      1317 ,    // 843
      1318 ,    // 844
      1320 ,    // 845
      1321 ,    // 846
      1323 ,    // 847
      1324 ,    // 848
      1326 ,    // 849
      1327 ,    // 850
      1329 ,    // 851
      1331 ,    // 852
      1332 ,    // 853
      1334 ,    // 854
      1335 ,    // 855
      1337 ,    // 856
      1338 ,    // 857
      1340 ,    // 858
      1341 ,    // 859
      1343 ,    // 860
      1345 ,    // 861
      1346 ,    // 862
      1348 ,    // 863
      1349 ,    // 864
      1351 ,    // 865
      1352 ,    // 866
      1354 ,    // 867
      1355 ,    // 868
      1357 ,    // 869
      1358 ,    // 870
      1360 ,    // 871
      1362 ,    // 872
      1363 ,    // 873
      1365 ,    // 874
      1366 ,    // 875
      1368 ,    // 876
      1369 ,    // 877
      1371 ,    // 878
      1372 ,    // 879
      1374 ,    // 880
      1375 ,    // 881
      1377 ,    // 882
      1379 ,    // 883
      1380 ,    // 884
      1382 ,    // 885
      1383 ,    // 886
      1385 ,    // 887
      1386 ,    // 888
      1388 ,    // 889
      1389 ,    // 890
      1391 ,    // 891
      1392 ,    // 892
      1394 ,    // 893
      1396 ,    // 894
      1397 ,    // 895
      1399 ,    // 896
      1400 ,    // 897
      1402 ,    // 898
      1403 ,    // 899
      1405 ,    // 900
      1406 ,    // 901
      1408 ,    // 902
      1409 ,    // 903
      1411 ,    // 904
      1413 ,    // 905
      1414 ,    // 906
      1416 ,    // 907
      1417 ,    // 908
      1419 ,    // 909
      1420 ,    // 910
      1422 ,    // 911
      1423 ,    // 912
      1425 ,    // 913
      1426 ,    // 914
      1428 ,    // 915
      1430 ,    // 916
      1431 ,    // 917
      1433 ,    // 918
      1434 ,    // 919
      1436 ,    // 920
      1437 ,    // 921
      1439 ,    // 922
      1440 ,    // 923
      1442 ,    // 924
      1443 ,    // 925
      1445 ,    // 926
      1447 ,    // 927
      1448 ,    // 928
      1450 ,    // 929
      1451 ,    // 930
      1453 ,    // 931
      1454 ,    // 932
      1456 ,    // 933
      1457 ,    // 934
      1459 ,    // 935
      1460 ,    // 936
      1462 ,    // 937
      1464 ,    // 938
      1465 ,    // 939
      1467 ,    // 940
      1468 ,    // 941
      1470 ,    // 942
      1471 ,    // 943
      1473 ,    // 944
      1474 ,    // 945
      1476 ,    // 946
      1477 ,    // 947
      1479 ,    // 948
      1480 ,    // 949
      1482 ,    // 950
      1484 ,    // 951
      1485 ,    // 952
      1487 ,    // 953
      1488 ,    // 954
      1490 ,    // 955
      1491 ,    // 956
      1493 ,    // 957
      1494 ,    // 958
      1496 ,    // 959
      1497 ,    // 960
      1499 ,    // 961
      1501 ,    // 962
      1502 ,    // 963
      1504 ,    // 964
      1505 ,    // 965
      1507 ,    // 966
      1508 ,    // 967
      1510 ,    // 968
      1511 ,    // 969
      1513 ,    // 970
      1514 ,    // 971
      1516 ,    // 972
      1518 ,    // 973
      1519 ,    // 974
      1521 ,    // 975
      1522 ,    // 976
      1524 ,    // 977
      1525 ,    // 978
      1527 ,    // 979
      1528 ,    // 980
      1530 ,    // 981
      1531 ,    // 982
      1533 ,    // 983
      1534 ,    // 984
      1536 ,    // 985
      1538 ,    // 986
      1539 ,    // 987
      1541 ,    // 988
      1542 ,    // 989
      1544 ,    // 990
      1545 ,    // 991
      1547 ,    // 992
      1548 ,    // 993
      1550 ,    // 994
      1551 ,    // 995
      1553 ,    // 996
      1554 ,    // 997
      1556 ,    // 998
      1558 ,    // 999
      1559 ,    // 1000
      1561 ,    // 1001
      1562 ,    // 1002
      1564 ,    // 1003
      1565 ,    // 1004
      1567 ,    // 1005
      1568 ,    // 1006
      1570 ,    // 1007
      1571 ,    // 1008
      1573 ,    // 1009
      1575 ,    // 1010
      1576 ,    // 1011
      1578 ,    // 1012
      1579 ,    // 1013
      1581 ,    // 1014
      1582 ,    // 1015
      1584 ,    // 1016
      1585 ,    // 1017
      1587 ,    // 1018
      1588 ,    // 1019
      1590 ,    // 1020
      1591 ,    // 1021
      1593 ,    // 1022
      1595 ,    // 1023
      1596 ,    // 1024
      1598 ,    // 1025
      1599 ,    // 1026
      1601 ,    // 1027
      1602 ,    // 1028
      1604 ,    // 1029
      1605 ,    // 1030
      1607 ,    // 1031
      1608 ,    // 1032
      1610 ,    // 1033
      1611 ,    // 1034
      1613 ,    // 1035
      1615 ,    // 1036
      1616 ,    // 1037
      1618 ,    // 1038
      1619 ,    // 1039
      1621 ,    // 1040
      1622 ,    // 1041
      1624 ,    // 1042
      1625 ,    // 1043
      1627 ,    // 1044
      1628 ,    // 1045
      1630 ,    // 1046
      1631 ,    // 1047
      1633 ,    // 1048
      1634 ,    // 1049
      1636 ,    // 1050
      1638 ,    // 1051
      1639 ,    // 1052
      1641 ,    // 1053
      1642 ,    // 1054
      1644 ,    // 1055
      1645 ,    // 1056
      1647 ,    // 1057
      1648 ,    // 1058
      1650 ,    // 1059
      1651 ,    // 1060
      1653 ,    // 1061
      1654 ,    // 1062
      1656 ,    // 1063
      1658 ,    // 1064
      1659 ,    // 1065
      1661 ,    // 1066
      1662 ,    // 1067
      1664 ,    // 1068
      1665 ,    // 1069
      1667 ,    // 1070
      1668 ,    // 1071
      1670 ,    // 1072
      1671 ,    // 1073
      1673 ,    // 1074
      1674 ,    // 1075
      1676 ,    // 1076
      1678 ,    // 1077
      1679 ,    // 1078
      1681 ,    // 1079
      1682 ,    // 1080
      1684 ,    // 1081
      1685 ,    // 1082
      1687 ,    // 1083
      1688 ,    // 1084
      1690 ,    // 1085
      1691 ,    // 1086
      1693 ,    // 1087
      1694 ,    // 1088
      1696 ,    // 1089
      1697 ,    // 1090
      1699 ,    // 1091
      1701 ,    // 1092
      1702 ,    // 1093
      1704 ,    // 1094
      1705 ,    // 1095
      1707 ,    // 1096
      1708 ,    // 1097
      1710 ,    // 1098
      1711 ,    // 1099
      1713 ,    // 1100
      1714 ,    // 1101
      1716 ,    // 1102
      1717 ,    // 1103
      1719 ,    // 1104
      1720 ,    // 1105
      1722 ,    // 1106
      1724 ,    // 1107
      1725 ,    // 1108
      1727 ,    // 1109
      1728 ,    // 1110
      1730 ,    // 1111
      1731 ,    // 1112
      1733 ,    // 1113
      1734 ,    // 1114
      1736 ,    // 1115
      1737 ,    // 1116
      1739 ,    // 1117
      1740 ,    // 1118
      1742 ,    // 1119
      1743 ,    // 1120
      1745 ,    // 1121
      1747 ,    // 1122
      1748 ,    // 1123
      1750 ,    // 1124
      1751 ,    // 1125
      1753 ,    // 1126
      1754 ,    // 1127
      1756 ,    // 1128
      1757 ,    // 1129
      1759 ,    // 1130
      1760 ,    // 1131
      1762 ,    // 1132
      1763 ,    // 1133
      1765 ,    // 1134
      1766 ,    // 1135
      1768 ,    // 1136
      1770 ,    // 1137
      1771 ,    // 1138
      1773 ,    // 1139
      1774 ,    // 1140
      1776 ,    // 1141
      1777 ,    // 1142
      1779 ,    // 1143
      1780 ,    // 1144
      1782 ,    // 1145
      1783 ,    // 1146
      1785 ,    // 1147
      1786 ,    // 1148
      1788 ,    // 1149
      1789 ,    // 1150
      1791 ,    // 1151
      1792 ,    // 1152
      1794 ,    // 1153
      1796 ,    // 1154
      1797 ,    // 1155
      1799 ,    // 1156
      1800 ,    // 1157
      1802 ,    // 1158
      1803 ,    // 1159
      1805 ,    // 1160
      1806 ,    // 1161
      1808 ,    // 1162
      1809 ,    // 1163
      1811 ,    // 1164
      1812 ,    // 1165
      1814 ,    // 1166
      1815 ,    // 1167
      1817 ,    // 1168
      1818 ,    // 1169
      1820 ,    // 1170
      1822 ,    // 1171
      1823 ,    // 1172
      1825 ,    // 1173
      1826 ,    // 1174
      1828 ,    // 1175
      1829 ,    // 1176
      1831 ,    // 1177
      1832 ,    // 1178
      1834 ,    // 1179
      1835 ,    // 1180
      1837 ,    // 1181
      1838 ,    // 1182
      1840 ,    // 1183
      1841 ,    // 1184
      1843 ,    // 1185
      1844 ,    // 1186
      1846 ,    // 1187
      1848 ,    // 1188
      1849 ,    // 1189
      1851 ,    // 1190
      1852 ,    // 1191
      1854 ,    // 1192
      1855 ,    // 1193
      1857 ,    // 1194
      1858 ,    // 1195
      1860 ,    // 1196
      1861 ,    // 1197
      1863 ,    // 1198
      1864 ,    // 1199
      1866 ,    // 1200
      1867 ,    // 1201
      1869 ,    // 1202
      1870 ,    // 1203
      1872 ,    // 1204
      1874 ,    // 1205
      1875 ,    // 1206
      1877 ,    // 1207
      1878 ,    // 1208
      1880 ,    // 1209
      1881 ,    // 1210
      1883 ,    // 1211
      1884 ,    // 1212
      1886 ,    // 1213
      1887 ,    // 1214
      1889 ,    // 1215
      1890 ,    // 1216
      1892 ,    // 1217
      1893 ,    // 1218
      1895 ,    // 1219
      1896 ,    // 1220
      1898 ,    // 1221
      1899 ,    // 1222
      1901 ,    // 1223
      1903 ,    // 1224
      1904 ,    // 1225
      1906 ,    // 1226
      1907 ,    // 1227
      1909 ,    // 1228
      1910 ,    // 1229
      1912 ,    // 1230
      1913 ,    // 1231
      1915 ,    // 1232
      1916 ,    // 1233
      1918 ,    // 1234
      1919 ,    // 1235
      1921 ,    // 1236
      1922 ,    // 1237
      1924 ,    // 1238
      1925 ,    // 1239
      1927 ,    // 1240
      1928 ,    // 1241
      1930 ,    // 1242
      1931 ,    // 1243
      1933 ,    // 1244
      1935 ,    // 1245
      1936 ,    // 1246
      1938 ,    // 1247
      1939 ,    // 1248
      1941 ,    // 1249
      1942 ,    // 1250
      1944 ,    // 1251
      1945 ,    // 1252
      1947 ,    // 1253
      1948 ,    // 1254
      1950 ,    // 1255
      1951 ,    // 1256
      1953 ,    // 1257
      1954 ,    // 1258
      1956 ,    // 1259
      1957 ,    // 1260
      1959 ,    // 1261
      1960 ,    // 1262
      1962 ,    // 1263
      1963 ,    // 1264
      1965 ,    // 1265
      1967 ,    // 1266
      1968 ,    // 1267
      1970 ,    // 1268
      1971 ,    // 1269
      1973 ,    // 1270
      1974 ,    // 1271
      1976 ,    // 1272
      1977 ,    // 1273
      1979 ,    // 1274
      1980 ,    // 1275
      1982 ,    // 1276
      1983 ,    // 1277
      1985 ,    // 1278
      1986 ,    // 1279
      1988 ,    // 1280
      1989 ,    // 1281
      1991 ,    // 1282
      1992 ,    // 1283
      1994 ,    // 1284
      1995 ,    // 1285
      1997 ,    // 1286
      1998 ,    // 1287
      2000 ,    // 1288
      2002 ,    // 1289
      2003 ,    // 1290
      2005 ,    // 1291
      2006 ,    // 1292
      2008 ,    // 1293
      2009 ,    // 1294
      2011 ,    // 1295
      2012 ,    // 1296
      2014 ,    // 1297
      2015 ,    // 1298
      2017 ,    // 1299
      2018 ,    // 1300
      2020 ,    // 1301
      2021 ,    // 1302
      2023 ,    // 1303
      2024 ,    // 1304
      2026 ,    // 1305
      2027 ,    // 1306
      2029 ,    // 1307
      2030 ,    // 1308
      2032 ,    // 1309
      2033 ,    // 1310
      2035 ,    // 1311
      2036 ,    // 1312
      2038 ,    // 1313
      2040 ,    // 1314
      2041 ,    // 1315
      2043 ,    // 1316
      2044 ,    // 1317
      2046 ,    // 1318
      2047 ,    // 1319
      2049 ,    // 1320
      2050 ,    // 1321
      2052 ,    // 1322
      2053 ,    // 1323
      2055 ,    // 1324
      2056 ,    // 1325
      2058 ,    // 1326
      2059 ,    // 1327
      2061 ,    // 1328
      2062 ,    // 1329
      2064 ,    // 1330
      2065 ,    // 1331
      2067 ,    // 1332
      2068 ,    // 1333
      2070 ,    // 1334
      2071 ,    // 1335
      2073 ,    // 1336
      2074 ,    // 1337
      2076 ,    // 1338
      2077 ,    // 1339
      2079 ,    // 1340
      2081 ,    // 1341
      2082 ,    // 1342
      2084 ,    // 1343
      2085 ,    // 1344
      2087 ,    // 1345
      2088 ,    // 1346
      2090 ,    // 1347
      2091 ,    // 1348
      2093 ,    // 1349
      2094 ,    // 1350
      2096 ,    // 1351
      2097 ,    // 1352
      2099 ,    // 1353
      2100 ,    // 1354
      2102 ,    // 1355
      2103 ,    // 1356
      2105 ,    // 1357
      2106 ,    // 1358
      2108 ,    // 1359
      2109 ,    // 1360
      2111 ,    // 1361
      2112 ,    // 1362
      2114 ,    // 1363
      2115 ,    // 1364
      2117 ,    // 1365
      2118 ,    // 1366
      2120 ,    // 1367
      2121 ,    // 1368
      2123 ,    // 1369
      2124 ,    // 1370
      2126 ,    // 1371
      2128 ,    // 1372
      2129 ,    // 1373
      2131 ,    // 1374
      2132 ,    // 1375
      2134 ,    // 1376
      2135 ,    // 1377
      2137 ,    // 1378
      2138 ,    // 1379
      2140 ,    // 1380
      2141 ,    // 1381
      2143 ,    // 1382
      2144 ,    // 1383
      2146 ,    // 1384
      2147 ,    // 1385
      2149 ,    // 1386
      2150 ,    // 1387
      2152 ,    // 1388
      2153 ,    // 1389
      2155 ,    // 1390
      2156 ,    // 1391
      2158 ,    // 1392
      2159 ,    // 1393
      2161 ,    // 1394
      2162 ,    // 1395
      2164 ,    // 1396
      2165 ,    // 1397
      2167 ,    // 1398
      2168 ,    // 1399
      2170 ,    // 1400
      2171 ,    // 1401
      2173 ,    // 1402
      2174 ,    // 1403
      2176 ,    // 1404
      2177 ,    // 1405
      2179 ,    // 1406
      2180 ,    // 1407
      2182 ,    // 1408
      2184 ,    // 1409
      2185 ,    // 1410
      2187 ,    // 1411
      2188 ,    // 1412
      2190 ,    // 1413
      2191 ,    // 1414
      2193 ,    // 1415
      2194 ,    // 1416
      2196 ,    // 1417
      2197 ,    // 1418
      2199 ,    // 1419
      2200 ,    // 1420
      2202 ,    // 1421
      2203 ,    // 1422
      2205 ,    // 1423
      2206 ,    // 1424
      2208 ,    // 1425
      2209 ,    // 1426
      2211 ,    // 1427
      2212 ,    // 1428
      2214 ,    // 1429
      2215 ,    // 1430
      2217 ,    // 1431
      2218 ,    // 1432
      2220 ,    // 1433
      2221 ,    // 1434
      2223 ,    // 1435
      2224 ,    // 1436
      2226 ,    // 1437
      2227 ,    // 1438
      2229 ,    // 1439
      2230 ,    // 1440
      2232 ,    // 1441
      2233 ,    // 1442
      2235 ,    // 1443
      2236 ,    // 1444
      2238 ,    // 1445
      2239 ,    // 1446
      2241 ,    // 1447
      2242 ,    // 1448
      2244 ,    // 1449
      2245 ,    // 1450
      2247 ,    // 1451
      2248 ,    // 1452
      2250 ,    // 1453
      2251 ,    // 1454
      2253 ,    // 1455
      2254 ,    // 1456
      2256 ,    // 1457
      2257 ,    // 1458
      2259 ,    // 1459
      2261 ,    // 1460
      2262 ,    // 1461
      2264 ,    // 1462
      2265 ,    // 1463
      2267 ,    // 1464
      2268 ,    // 1465
      2270 ,    // 1466
      2271 ,    // 1467
      2273 ,    // 1468
      2274 ,    // 1469
      2276 ,    // 1470
      2277 ,    // 1471
      2279 ,    // 1472
      2280 ,    // 1473
      2282 ,    // 1474
      2283 ,    // 1475
      2285 ,    // 1476
      2286 ,    // 1477
      2288 ,    // 1478
      2289 ,    // 1479
      2291 ,    // 1480
      2292 ,    // 1481
      2294 ,    // 1482
      2295 ,    // 1483
      2297 ,    // 1484
      2298 ,    // 1485
      2300 ,    // 1486
      2301 ,    // 1487
      2303 ,    // 1488
      2304 ,    // 1489
      2306 ,    // 1490
      2307 ,    // 1491
      2309 ,    // 1492
      2310 ,    // 1493
      2312 ,    // 1494
      2313 ,    // 1495
      2315 ,    // 1496
      2316 ,    // 1497
      2318 ,    // 1498
      2319 ,    // 1499
      2321 ,    // 1500
      2322 ,    // 1501
      2324 ,    // 1502
      2325 ,    // 1503
      2327 ,    // 1504
      2328 ,    // 1505
      2330 ,    // 1506
      2331 ,    // 1507
      2333 ,    // 1508
      2334 ,    // 1509
      2336 ,    // 1510
      2337 ,    // 1511
      2339 ,    // 1512
      2340 ,    // 1513
      2342 ,    // 1514
      2343 ,    // 1515
      2345 ,    // 1516
      2346 ,    // 1517
      2348 ,    // 1518
      2349 ,    // 1519
      2351 ,    // 1520
      2352 ,    // 1521
      2354 ,    // 1522
      2355 ,    // 1523
      2357 ,    // 1524
      2358 ,    // 1525
      2360 ,    // 1526
      2361 ,    // 1527
      2363 ,    // 1528
      2364 ,    // 1529
      2366 ,    // 1530
      2367 ,    // 1531
      2369 ,    // 1532
      2370 ,    // 1533
      2372 ,    // 1534
      2373 ,    // 1535
      2375 ,    // 1536
      2376 ,    // 1537
      2378 ,    // 1538
      2379 ,    // 1539
      2381 ,    // 1540
      2382 ,    // 1541
      2384 ,    // 1542
      2385 ,    // 1543
      2387 ,    // 1544
      2388 ,    // 1545
      2390 ,    // 1546
      2391 ,    // 1547
      2393 ,    // 1548
      2394 ,    // 1549
      2396 ,    // 1550
      2397 ,    // 1551
      2399 ,    // 1552
      2400 ,    // 1553
      2402 ,    // 1554
      2403 ,    // 1555
      2405 ,    // 1556
      2406 ,    // 1557
      2408 ,    // 1558
      2409 ,    // 1559
      2411 ,    // 1560
      2412 ,    // 1561
      2414 ,    // 1562
      2415 ,    // 1563
      2417 ,    // 1564
      2418 ,    // 1565
      2420 ,    // 1566
      2421 ,    // 1567
      2423 ,    // 1568
      2424 ,    // 1569
      2426 ,    // 1570
      2427 ,    // 1571
      2429 ,    // 1572
      2430 ,    // 1573
      2432 ,    // 1574
      2433 ,    // 1575
      2435 ,    // 1576
      2436 ,    // 1577
      2438 ,    // 1578
      2439 ,    // 1579
      2441 ,    // 1580
      2442 ,    // 1581
      2444 ,    // 1582
      2445 ,    // 1583
      2447 ,    // 1584
      2448 ,    // 1585
      2450 ,    // 1586
      2451 ,    // 1587
      2453 ,    // 1588
      2454 ,    // 1589
      2456 ,    // 1590
      2457 ,    // 1591
      2459 ,    // 1592
      2460 ,    // 1593
      2462 ,    // 1594
      2463 ,    // 1595
      2465 ,    // 1596
      2466 ,    // 1597
      2468 ,    // 1598
      2469 ,    // 1599
      2471 ,    // 1600
      2472 ,    // 1601
      2474 ,    // 1602
      2475 ,    // 1603
      2477 ,    // 1604
      2478 ,    // 1605
      2480 ,    // 1606
      2481 ,    // 1607
      2483 ,    // 1608
      2484 ,    // 1609
      2486 ,    // 1610
      2487 ,    // 1611
      2489 ,    // 1612
      2490 ,    // 1613
      2492 ,    // 1614
      2493 ,    // 1615
      2495 ,    // 1616
      2496 ,    // 1617
      2498 ,    // 1618
      2499 ,    // 1619
      2501 ,    // 1620
      2502 ,    // 1621
      2504 ,    // 1622
      2505 ,    // 1623
      2507 ,    // 1624
      2508 ,    // 1625
      2510 ,    // 1626
      2511 ,    // 1627
      2513 ,    // 1628
      2514 ,    // 1629
      2516 ,    // 1630
      2517 ,    // 1631
      2519 ,    // 1632
      2520 ,    // 1633
      2522 ,    // 1634
      2523 ,    // 1635
      2525 ,    // 1636
      2526 ,    // 1637
      2527 ,    // 1638
      2529 ,    // 1639
      2530 ,    // 1640
      2532 ,    // 1641
      2533 ,    // 1642
      2535 ,    // 1643
      2536 ,    // 1644
      2538 ,    // 1645
      2539 ,    // 1646
      2541 ,    // 1647
      2542 ,    // 1648
      2544 ,    // 1649
      2545 ,    // 1650
      2547 ,    // 1651
      2548 ,    // 1652
      2550 ,    // 1653
      2551 ,    // 1654
      2553 ,    // 1655
      2554 ,    // 1656
      2556 ,    // 1657
      2557 ,    // 1658
      2559 ,    // 1659
      2560 ,    // 1660
      2562 ,    // 1661
      2563 ,    // 1662
      2565 ,    // 1663
      2566 ,    // 1664
      2568 ,    // 1665
      2569 ,    // 1666
      2571 ,    // 1667
      2572 ,    // 1668
      2574 ,    // 1669
      2575 ,    // 1670
      2577 ,    // 1671
      2578 ,    // 1672
      2580 ,    // 1673
      2581 ,    // 1674
      2583 ,    // 1675
      2584 ,    // 1676
      2586 ,    // 1677
      2587 ,    // 1678
      2589 ,    // 1679
      2590 ,    // 1680
      2592 ,    // 1681
      2593 ,    // 1682
      2595 ,    // 1683
      2596 ,    // 1684
      2598 ,    // 1685
      2599 ,    // 1686
      2600 ,    // 1687
      2602 ,    // 1688
      2603 ,    // 1689
      2605 ,    // 1690
      2606 ,    // 1691
      2608 ,    // 1692
      2609 ,    // 1693
      2611 ,    // 1694
      2612 ,    // 1695
      2614 ,    // 1696
      2615 ,    // 1697
      2617 ,    // 1698
      2618 ,    // 1699
      2620 ,    // 1700
      2621 ,    // 1701
      2623 ,    // 1702
      2624 ,    // 1703
      2626 ,    // 1704
      2627 ,    // 1705
      2629 ,    // 1706
      2630 ,    // 1707
      2632 ,    // 1708
      2633 ,    // 1709
      2635 ,    // 1710
      2636 ,    // 1711
      2638 ,    // 1712
      2639 ,    // 1713
      2641 ,    // 1714
      2642 ,    // 1715
      2644 ,    // 1716
      2645 ,    // 1717
      2647 ,    // 1718
      2648 ,    // 1719
      2650 ,    // 1720
      2651 ,    // 1721
      2652 ,    // 1722
      2654 ,    // 1723
      2655 ,    // 1724
      2657 ,    // 1725
      2658 ,    // 1726
      2660 ,    // 1727
      2661 ,    // 1728
      2663 ,    // 1729
      2664 ,    // 1730
      2666 ,    // 1731
      2667 ,    // 1732
      2669 ,    // 1733
      2670 ,    // 1734
      2672 ,    // 1735
      2673 ,    // 1736
      2675 ,    // 1737
      2676 ,    // 1738
      2678 ,    // 1739
      2679 ,    // 1740
      2681 ,    // 1741
      2682 ,    // 1742
      2684 ,    // 1743
      2685 ,    // 1744
      2687 ,    // 1745
      2688 ,    // 1746
      2690 ,    // 1747
      2691 ,    // 1748
      2693 ,    // 1749
      2694 ,    // 1750
      2695 ,    // 1751
      2697 ,    // 1752
      2698 ,    // 1753
      2700 ,    // 1754
      2701 ,    // 1755
      2703 ,    // 1756
      2704 ,    // 1757
      2706 ,    // 1758
      2707 ,    // 1759
      2709 ,    // 1760
      2710 ,    // 1761
      2712 ,    // 1762
      2713 ,    // 1763
      2715 ,    // 1764
      2716 ,    // 1765
      2718 ,    // 1766
      2719 ,    // 1767
      2721 ,    // 1768
      2722 ,    // 1769
      2724 ,    // 1770
      2725 ,    // 1771
      2727 ,    // 1772
      2728 ,    // 1773
      2730 ,    // 1774
      2731 ,    // 1775
      2732 ,    // 1776
      2734 ,    // 1777
      2735 ,    // 1778
      2737 ,    // 1779
      2738 ,    // 1780
      2740 ,    // 1781
      2741 ,    // 1782
      2743 ,    // 1783
      2744 ,    // 1784
      2746 ,    // 1785
      2747 ,    // 1786
      2749 ,    // 1787
      2750 ,    // 1788
      2752 ,    // 1789
      2753 ,    // 1790
      2755 ,    // 1791
      2756 ,    // 1792
      2758 ,    // 1793
      2759 ,    // 1794
      2761 ,    // 1795
      2762 ,    // 1796
      2764 ,    // 1797
      2765 ,    // 1798
      2766 ,    // 1799
      2768 ,    // 1800
      2769 ,    // 1801
      2771 ,    // 1802
      2772 ,    // 1803
      2774 ,    // 1804
      2775 ,    // 1805
      2777 ,    // 1806
      2778 ,    // 1807
      2780 ,    // 1808
      2781 ,    // 1809
      2783 ,    // 1810
      2784 ,    // 1811
      2786 ,    // 1812
      2787 ,    // 1813
      2789 ,    // 1814
      2790 ,    // 1815
      2792 ,    // 1816
      2793 ,    // 1817
      2794 ,    // 1818
      2796 ,    // 1819
      2797 ,    // 1820
      2799 ,    // 1821
      2800 ,    // 1822
      2802 ,    // 1823
      2803 ,    // 1824
      2805 ,    // 1825
      2806 ,    // 1826
      2808 ,    // 1827
      2809 ,    // 1828
      2811 ,    // 1829
      2812 ,    // 1830
      2814 ,    // 1831
      2815 ,    // 1832
      2817 ,    // 1833
      2818 ,    // 1834
      2820 ,    // 1835
      2821 ,    // 1836
      2822 ,    // 1837
      2824 ,    // 1838
      2825 ,    // 1839
      2827 ,    // 1840
      2828 ,    // 1841
      2830 ,    // 1842
      2831 ,    // 1843
      2833 ,    // 1844
      2834 ,    // 1845
      2836 ,    // 1846
      2837 ,    // 1847
      2839 ,    // 1848
      2840 ,    // 1849
      2842 ,    // 1850
      2843 ,    // 1851
      2845 ,    // 1852
      2846 ,    // 1853
      2847 ,    // 1854
      2849 ,    // 1855
      2850 ,    // 1856
      2852 ,    // 1857
      2853 ,    // 1858
      2855 ,    // 1859
      2856 ,    // 1860
      2858 ,    // 1861
      2859 ,    // 1862
      2861 ,    // 1863
      2862 ,    // 1864
      2864 ,    // 1865
      2865 ,    // 1866
      2867 ,    // 1867
      2868 ,    // 1868
      2870 ,    // 1869
      2871 ,    // 1870
      2872 ,    // 1871
      2874 ,    // 1872
      2875 ,    // 1873
      2877 ,    // 1874
      2878 ,    // 1875
      2880 ,    // 1876
      2881 ,    // 1877
      2883 ,    // 1878
      2884 ,    // 1879
      2886 ,    // 1880
      2887 ,    // 1881
      2889 ,    // 1882
      2890 ,    // 1883
      2892 ,    // 1884
      2893 ,    // 1885
      2894 ,    // 1886
      2896 ,    // 1887
      2897 ,    // 1888
      2899 ,    // 1889
      2900 ,    // 1890
      2902 ,    // 1891
      2903 ,    // 1892
      2905 ,    // 1893
      2906 ,    // 1894
      2908 ,    // 1895
      2909 ,    // 1896
      2911 ,    // 1897
      2912 ,    // 1898
      2914 ,    // 1899
      2915 ,    // 1900
      2916 ,    // 1901
      2918 ,    // 1902
      2919 ,    // 1903
      2921 ,    // 1904
      2922 ,    // 1905
      2924 ,    // 1906
      2925 ,    // 1907
      2927 ,    // 1908
      2928 ,    // 1909
      2930 ,    // 1910
      2931 ,    // 1911
      2933 ,    // 1912
      2934 ,    // 1913
      2936 ,    // 1914
      2937 ,    // 1915
      2938 ,    // 1916
      2940 ,    // 1917
      2941 ,    // 1918
      2943 ,    // 1919
      2944 ,    // 1920
      2946 ,    // 1921
      2947 ,    // 1922
      2949 ,    // 1923
      2950 ,    // 1924
      2952 ,    // 1925
      2953 ,    // 1926
      2955 ,    // 1927
      2956 ,    // 1928
      2957 ,    // 1929
      2959 ,    // 1930
      2960 ,    // 1931
      2962 ,    // 1932
      2963 ,    // 1933
      2965 ,    // 1934
      2966 ,    // 1935
      2968 ,    // 1936
      2969 ,    // 1937
      2971 ,    // 1938
      2972 ,    // 1939
      2974 ,    // 1940
      2975 ,    // 1941
      2976 ,    // 1942
      2978 ,    // 1943
      2979 ,    // 1944
      2981 ,    // 1945
      2982 ,    // 1946
      2984 ,    // 1947
      2985 ,    // 1948
      2987 ,    // 1949
      2988 ,    // 1950
      2990 ,    // 1951
      2991 ,    // 1952
      2993 ,    // 1953
      2994 ,    // 1954
      2995 ,    // 1955
      2997 ,    // 1956
      2998 ,    // 1957
      3000 ,    // 1958
      3001 ,    // 1959
      3003 ,    // 1960
      3004 ,    // 1961
      3006 ,    // 1962
      3007 ,    // 1963
      3009 ,    // 1964
      3010 ,    // 1965
      3012 ,    // 1966
      3013 ,    // 1967
      3014 ,    // 1968
      3016 ,    // 1969
      3017 ,    // 1970
      3019 ,    // 1971
      3020 ,    // 1972
      3022 ,    // 1973
      3023 ,    // 1974
      3025 ,    // 1975
      3026 ,    // 1976
      3028 ,    // 1977
      3029 ,    // 1978
      3030 ,    // 1979
      3032 ,    // 1980
      3033 ,    // 1981
      3035 ,    // 1982
      3036 ,    // 1983
      3038 ,    // 1984
      3039 ,    // 1985
      3041 ,    // 1986
      3042 ,    // 1987
      3044 ,    // 1988
      3045 ,    // 1989
      3047 ,    // 1990
      3048 ,    // 1991
      3049 ,    // 1992
      3051 ,    // 1993
      3052 ,    // 1994
      3054 ,    // 1995
      3055 ,    // 1996
      3057 ,    // 1997
      3058 ,    // 1998
      3060 ,    // 1999
      3061 ,    // 2000
      3063 ,    // 2001
      3064 ,    // 2002
      3065 ,    // 2003
      3067 ,    // 2004
      3068 ,    // 2005
      3070 ,    // 2006
      3071 ,    // 2007
      3073 ,    // 2008
      3074 ,    // 2009
      3076 ,    // 2010
      3077 ,    // 2011
      3079 ,    // 2012
      3080 ,    // 2013
      3081 ,    // 2014
      3083 ,    // 2015
      3084 ,    // 2016
      3086 ,    // 2017
      3087 ,    // 2018
      3089 ,    // 2019
      3090 ,    // 2020
      3092 ,    // 2021
      3093 ,    // 2022
      3094 ,    // 2023
      3096 ,    // 2024
      3097 ,    // 2025
      3099 ,    // 2026
      3100 ,    // 2027
      3102 ,    // 2028
      3103 ,    // 2029
      3105 ,    // 2030
      3106 ,    // 2031
      3108 ,    // 2032
      3109 ,    // 2033
      3110 ,    // 2034
      3112 ,    // 2035
      3113 ,    // 2036
      3115 ,    // 2037
      3116 ,    // 2038
      3118 ,    // 2039
      3119 ,    // 2040
      3121 ,    // 2041
      3122 ,    // 2042
      3124 ,    // 2043
      3125 ,    // 2044
      3126 ,    // 2045
      3128 ,    // 2046
      3129 ,    // 2047
      3131 ,    // 2048
      3132 ,    // 2049
      3134 ,    // 2050
      3135 ,    // 2051
      3137 ,    // 2052
      3138 ,    // 2053
      3139 ,    // 2054
      3141 ,    // 2055
      3142 ,    // 2056
      3144 ,    // 2057
      3145 ,    // 2058
      3147 ,    // 2059
      3148 ,    // 2060
      3150 ,    // 2061
      3151 ,    // 2062
      3152 ,    // 2063
      3154 ,    // 2064
      3155 ,    // 2065
      3157 ,    // 2066
      3158 ,    // 2067
      3160 ,    // 2068
      3161 ,    // 2069
      3163 ,    // 2070
      3164 ,    // 2071
      3166 ,    // 2072
      3167 ,    // 2073
      3168 ,    // 2074
      3170 ,    // 2075
      3171 ,    // 2076
      3173 ,    // 2077
      3174 ,    // 2078
      3176 ,    // 2079
      3177 ,    // 2080
      3179 ,    // 2081
      3180 ,    // 2082
      3181 ,    // 2083
      3183 ,    // 2084
      3184 ,    // 2085
      3186 ,    // 2086
      3187 ,    // 2087
      3189 ,    // 2088
      3190 ,    // 2089
      3192 ,    // 2090
      3193 ,    // 2091
      3194 ,    // 2092
      3196 ,    // 2093
      3197 ,    // 2094
      3199 ,    // 2095
      3200 ,    // 2096
      3202 ,    // 2097
      3203 ,    // 2098
      3205 ,    // 2099
      3206 ,    // 2100
      3207 ,    // 2101
      3209 ,    // 2102
      3210 ,    // 2103
      3212 ,    // 2104
      3213 ,    // 2105
      3215 ,    // 2106
      3216 ,    // 2107
      3218 ,    // 2108
      3219 ,    // 2109
      3220 ,    // 2110
      3222 ,    // 2111
      3223 ,    // 2112
      3225 ,    // 2113
      3226 ,    // 2114
      3228 ,    // 2115
      3229 ,    // 2116
      3230 ,    // 2117
      3232 ,    // 2118
      3233 ,    // 2119
      3235 ,    // 2120
      3236 ,    // 2121
      3238 ,    // 2122
      3239 ,    // 2123
      3241 ,    // 2124
      3242 ,    // 2125
      3243 ,    // 2126
      3245 ,    // 2127
      3246 ,    // 2128
      3248 ,    // 2129
      3249 ,    // 2130
      3251 ,    // 2131
      3252 ,    // 2132
      3254 ,    // 2133
      3255 ,    // 2134
      3256 ,    // 2135
      3258 ,    // 2136
      3259 ,    // 2137
      3261 ,    // 2138
      3262 ,    // 2139
      3264 ,    // 2140
      3265 ,    // 2141
      3266 ,    // 2142
      3268 ,    // 2143
      3269 ,    // 2144
      3271 ,    // 2145
      3272 ,    // 2146
      3274 ,    // 2147
      3275 ,    // 2148
      3277 ,    // 2149
      3278 ,    // 2150
      3279 ,    // 2151
      3281 ,    // 2152
      3282 ,    // 2153
      3284 ,    // 2154
      3285 ,    // 2155
      3287 ,    // 2156
      3288 ,    // 2157
      3289 ,    // 2158
      3291 ,    // 2159
      3292 ,    // 2160
      3294 ,    // 2161
      3295 ,    // 2162
      3297 ,    // 2163
      3298 ,    // 2164
      3300 ,    // 2165
      3301 ,    // 2166
      3302 ,    // 2167
      3304 ,    // 2168
      3305 ,    // 2169
      3307 ,    // 2170
      3308 ,    // 2171
      3310 ,    // 2172
      3311 ,    // 2173
      3312 ,    // 2174
      3314 ,    // 2175
      3315 ,    // 2176
      3317 ,    // 2177
      3318 ,    // 2178
      3320 ,    // 2179
      3321 ,    // 2180
      3322 ,    // 2181
      3324 ,    // 2182
      3325 ,    // 2183
      3327 ,    // 2184
      3328 ,    // 2185
      3330 ,    // 2186
      3331 ,    // 2187
      3333 ,    // 2188
      3334 ,    // 2189
      3335 ,    // 2190
      3337 ,    // 2191
      3338 ,    // 2192
      3340 ,    // 2193
      3341 ,    // 2194
      3343 ,    // 2195
      3344 ,    // 2196
      3345 ,    // 2197
      3347 ,    // 2198
      3348 ,    // 2199
      3350 ,    // 2200
      3351 ,    // 2201
      3353 ,    // 2202
      3354 ,    // 2203
      3355 ,    // 2204
      3357 ,    // 2205
      3358 ,    // 2206
      3360 ,    // 2207
      3361 ,    // 2208
      3363 ,    // 2209
      3364 ,    // 2210
      3365 ,    // 2211
      3367 ,    // 2212
      3368 ,    // 2213
      3370 ,    // 2214
      3371 ,    // 2215
      3373 ,    // 2216
      3374 ,    // 2217
      3375 ,    // 2218
      3377 ,    // 2219
      3378 ,    // 2220
      3380 ,    // 2221
      3381 ,    // 2222
      3383 ,    // 2223
      3384 ,    // 2224
      3385 ,    // 2225
      3387 ,    // 2226
      3388 ,    // 2227
      3390 ,    // 2228
      3391 ,    // 2229
      3393 ,    // 2230
      3394 ,    // 2231
      3395 ,    // 2232
      3397 ,    // 2233
      3398 ,    // 2234
      3400 ,    // 2235
      3401 ,    // 2236
      3403 ,    // 2237
      3404 ,    // 2238
      3405 ,    // 2239
      3407 ,    // 2240
      3408 ,    // 2241
      3410 ,    // 2242
      3411 ,    // 2243
      3413 ,    // 2244
      3414 ,    // 2245
      3415 ,    // 2246
      3417 ,    // 2247
      3418 ,    // 2248
      3420 ,    // 2249
      3421 ,    // 2250
      3423 ,    // 2251
      3424 ,    // 2252
      3425 ,    // 2253
      3427 ,    // 2254
      3428 ,    // 2255
      3430 ,    // 2256
      3431 ,    // 2257
      3432 ,    // 2258
      3434 ,    // 2259
      3435 ,    // 2260
      3437 ,    // 2261
      3438 ,    // 2262
      3440 ,    // 2263
      3441 ,    // 2264
      3442 ,    // 2265
      3444 ,    // 2266
      3445 ,    // 2267
      3447 ,    // 2268
      3448 ,    // 2269
      3450 ,    // 2270
      3451 ,    // 2271
      3452 ,    // 2272
      3454 ,    // 2273
      3455 ,    // 2274
      3457 ,    // 2275
      3458 ,    // 2276
      3460 ,    // 2277
      3461 ,    // 2278
      3462 ,    // 2279
      3464 ,    // 2280
      3465 ,    // 2281
      3467 ,    // 2282
      3468 ,    // 2283
      3469 ,    // 2284
      3471 ,    // 2285
      3472 ,    // 2286
      3474 ,    // 2287
      3475 ,    // 2288
      3477 ,    // 2289
      3478 ,    // 2290
      3479 ,    // 2291
      3481 ,    // 2292
      3482 ,    // 2293
      3484 ,    // 2294
      3485 ,    // 2295
      3487 ,    // 2296
      3488 ,    // 2297
      3489 ,    // 2298
      3491 ,    // 2299
      3492 ,    // 2300
      3494 ,    // 2301
      3495 ,    // 2302
      3496 ,    // 2303
      3498 ,    // 2304
      3499 ,    // 2305
      3501 ,    // 2306
      3502 ,    // 2307
      3504 ,    // 2308
      3505 ,    // 2309
      3506 ,    // 2310
      3508 ,    // 2311
      3509 ,    // 2312
      3511 ,    // 2313
      3512 ,    // 2314
      3513 ,    // 2315
      3515 ,    // 2316
      3516 ,    // 2317
      3518 ,    // 2318
      3519 ,    // 2319
      3521 ,    // 2320
      3522 ,    // 2321
      3523 ,    // 2322
      3525 ,    // 2323
      3526 ,    // 2324
      3528 ,    // 2325
      3529 ,    // 2326
      3530 ,    // 2327
      3532 ,    // 2328
      3533 ,    // 2329
      3535 ,    // 2330
      3536 ,    // 2331
      3538 ,    // 2332
      3539 ,    // 2333
      3540 ,    // 2334
      3542 ,    // 2335
      3543 ,    // 2336
      3545 ,    // 2337
      3546 ,    // 2338
      3547 ,    // 2339
      3549 ,    // 2340
      3550 ,    // 2341
      3552 ,    // 2342
      3553 ,    // 2343
      3554 ,    // 2344
      3556 ,    // 2345
      3557 ,    // 2346
      3559 ,    // 2347
      3560 ,    // 2348
      3562 ,    // 2349
      3563 ,    // 2350
      3564 ,    // 2351
      3566 ,    // 2352
      3567 ,    // 2353
      3569 ,    // 2354
      3570 ,    // 2355
      3571 ,    // 2356
      3573 ,    // 2357
      3574 ,    // 2358
      3576 ,    // 2359
      3577 ,    // 2360
      3578 ,    // 2361
      3580 ,    // 2362
      3581 ,    // 2363
      3583 ,    // 2364
      3584 ,    // 2365
      3586 ,    // 2366
      3587 ,    // 2367
      3588 ,    // 2368
      3590 ,    // 2369
      3591 ,    // 2370
      3593 ,    // 2371
      3594 ,    // 2372
      3595 ,    // 2373
      3597 ,    // 2374
      3598 ,    // 2375
      3600 ,    // 2376
      3601 ,    // 2377
      3602 ,    // 2378
      3604 ,    // 2379
      3605 ,    // 2380
      3607 ,    // 2381
      3608 ,    // 2382
      3609 ,    // 2383
      3611 ,    // 2384
      3612 ,    // 2385
      3614 ,    // 2386
      3615 ,    // 2387
      3617 ,    // 2388
      3618 ,    // 2389
      3619 ,    // 2390
      3621 ,    // 2391
      3622 ,    // 2392
      3624 ,    // 2393
      3625 ,    // 2394
      3626 ,    // 2395
      3628 ,    // 2396
      3629 ,    // 2397
      3631 ,    // 2398
      3632 ,    // 2399
      3633 ,    // 2400
      3635 ,    // 2401
      3636 ,    // 2402
      3638 ,    // 2403
      3639 ,    // 2404
      3640 ,    // 2405
      3642 ,    // 2406
      3643 ,    // 2407
      3645 ,    // 2408
      3646 ,    // 2409
      3647 ,    // 2410
      3649 ,    // 2411
      3650 ,    // 2412
      3652 ,    // 2413
      3653 ,    // 2414
      3654 ,    // 2415
      3656 ,    // 2416
      3657 ,    // 2417
      3659 ,    // 2418
      3660 ,    // 2419
      3661 ,    // 2420
      3663 ,    // 2421
      3664 ,    // 2422
      3666 ,    // 2423
      3667 ,    // 2424
      3668 ,    // 2425
      3670 ,    // 2426
      3671 ,    // 2427
      3673 ,    // 2428
      3674 ,    // 2429
      3675 ,    // 2430
      3677 ,    // 2431
      3678 ,    // 2432
      3680 ,    // 2433
      3681 ,    // 2434
      3683 ,    // 2435
      3684 ,    // 2436
      3685 ,    // 2437
      3687 ,    // 2438
      3688 ,    // 2439
      3690 ,    // 2440
      3691 ,    // 2441
      3692 ,    // 2442
      3694 ,    // 2443
      3695 ,    // 2444
      3697 ,    // 2445
      3698 ,    // 2446
      3699 ,    // 2447
      3701 ,    // 2448
      3702 ,    // 2449
      3703 ,    // 2450
      3705 ,    // 2451
      3706 ,    // 2452
      3708 ,    // 2453
      3709 ,    // 2454
      3710 ,    // 2455
      3712 ,    // 2456
      3713 ,    // 2457
      3715 ,    // 2458
      3716 ,    // 2459
      3717 ,    // 2460
      3719 ,    // 2461
      3720 ,    // 2462
      3722 ,    // 2463
      3723 ,    // 2464
      3724 ,    // 2465
      3726 ,    // 2466
      3727 ,    // 2467
      3729 ,    // 2468
      3730 ,    // 2469
      3731 ,    // 2470
      3733 ,    // 2471
      3734 ,    // 2472
      3736 ,    // 2473
      3737 ,    // 2474
      3738 ,    // 2475
      3740 ,    // 2476
      3741 ,    // 2477
      3743 ,    // 2478
      3744 ,    // 2479
      3745 ,    // 2480
      3747 ,    // 2481
      3748 ,    // 2482
      3750 ,    // 2483
      3751 ,    // 2484
      3752 ,    // 2485
      3754 ,    // 2486
      3755 ,    // 2487
      3757 ,    // 2488
      3758 ,    // 2489
      3759 ,    // 2490
      3761 ,    // 2491
      3762 ,    // 2492
      3764 ,    // 2493
      3765 ,    // 2494
      3766 ,    // 2495
      3768 ,    // 2496
      3769 ,    // 2497
      3770 ,    // 2498
      3772 ,    // 2499
      3773 ,    // 2500
      3775 ,    // 2501
      3776 ,    // 2502
      3777 ,    // 2503
      3779 ,    // 2504
      3780 ,    // 2505
      3782 ,    // 2506
      3783 ,    // 2507
      3784 ,    // 2508
      3786 ,    // 2509
      3787 ,    // 2510
      3789 ,    // 2511
      3790 ,    // 2512
      3791 ,    // 2513
      3793 ,    // 2514
      3794 ,    // 2515
      3796 ,    // 2516
      3797 ,    // 2517
      3798 ,    // 2518
      3800 ,    // 2519
      3801 ,    // 2520
      3802 ,    // 2521
      3804 ,    // 2522
      3805 ,    // 2523
      3807 ,    // 2524
      3808 ,    // 2525
      3809 ,    // 2526
      3811 ,    // 2527
      3812 ,    // 2528
      3814 ,    // 2529
      3815 ,    // 2530
      3816 ,    // 2531
      3818 ,    // 2532
      3819 ,    // 2533
      3821 ,    // 2534
      3822 ,    // 2535
      3823 ,    // 2536
      3825 ,    // 2537
      3826 ,    // 2538
      3827 ,    // 2539
      3829 ,    // 2540
      3830 ,    // 2541
      3832 ,    // 2542
      3833 ,    // 2543
      3834 ,    // 2544
      3836 ,    // 2545
      3837 ,    // 2546
      3839 ,    // 2547
      3840 ,    // 2548
      3841 ,    // 2549
      3843 ,    // 2550
      3844 ,    // 2551
      3845 ,    // 2552
      3847 ,    // 2553
      3848 ,    // 2554
      3850 ,    // 2555
      3851 ,    // 2556
      3852 ,    // 2557
      3854 ,    // 2558
      3855 ,    // 2559
      3857 ,    // 2560
      3858 ,    // 2561
      3859 ,    // 2562
      3861 ,    // 2563
      3862 ,    // 2564
      3863 ,    // 2565
      3865 ,    // 2566
      3866 ,    // 2567
      3868 ,    // 2568
      3869 ,    // 2569
      3870 ,    // 2570
      3872 ,    // 2571
      3873 ,    // 2572
      3874 ,    // 2573
      3876 ,    // 2574
      3877 ,    // 2575
      3879 ,    // 2576
      3880 ,    // 2577
      3881 ,    // 2578
      3883 ,    // 2579
      3884 ,    // 2580
      3886 ,    // 2581
      3887 ,    // 2582
      3888 ,    // 2583
      3890 ,    // 2584
      3891 ,    // 2585
      3892 ,    // 2586
      3894 ,    // 2587
      3895 ,    // 2588
      3897 ,    // 2589
      3898 ,    // 2590
      3899 ,    // 2591
      3901 ,    // 2592
      3902 ,    // 2593
      3903 ,    // 2594
      3905 ,    // 2595
      3906 ,    // 2596
      3908 ,    // 2597
      3909 ,    // 2598
      3910 ,    // 2599
      3912 ,    // 2600
      3913 ,    // 2601
      3915 ,    // 2602
      3916 ,    // 2603
      3917 ,    // 2604
      3919 ,    // 2605
      3920 ,    // 2606
      3921 ,    // 2607
      3923 ,    // 2608
      3924 ,    // 2609
      3926 ,    // 2610
      3927 ,    // 2611
      3928 ,    // 2612
      3930 ,    // 2613
      3931 ,    // 2614
      3932 ,    // 2615
      3934 ,    // 2616
      3935 ,    // 2617
      3937 ,    // 2618
      3938 ,    // 2619
      3939 ,    // 2620
      3941 ,    // 2621
      3942 ,    // 2622
      3943 ,    // 2623
      3945 ,    // 2624
      3946 ,    // 2625
      3948 ,    // 2626
      3949 ,    // 2627
      3950 ,    // 2628
      3952 ,    // 2629
      3953 ,    // 2630
      3954 ,    // 2631
      3956 ,    // 2632
      3957 ,    // 2633
      3959 ,    // 2634
      3960 ,    // 2635
      3961 ,    // 2636
      3963 ,    // 2637
      3964 ,    // 2638
      3965 ,    // 2639
      3967 ,    // 2640
      3968 ,    // 2641
      3969 ,    // 2642
      3971 ,    // 2643
      3972 ,    // 2644
      3974 ,    // 2645
      3975 ,    // 2646
      3976 ,    // 2647
      3978 ,    // 2648
      3979 ,    // 2649
      3980 ,    // 2650
      3982 ,    // 2651
      3983 ,    // 2652
      3985 ,    // 2653
      3986 ,    // 2654
      3987 ,    // 2655
      3989 ,    // 2656
      3990 ,    // 2657
      3991 ,    // 2658
      3993 ,    // 2659
      3994 ,    // 2660
      3996 ,    // 2661
      3997 ,    // 2662
      3998 ,    // 2663
      4000 ,    // 2664
      4001 ,    // 2665
      4002 ,    // 2666
      4004 ,    // 2667
      4005 ,    // 2668
      4006 ,    // 2669
      4008 ,    // 2670
      4009 ,    // 2671
      4011 ,    // 2672
      4012 ,    // 2673
      4013 ,    // 2674
      4015 ,    // 2675
      4016 ,    // 2676
      4017 ,    // 2677
      4019 ,    // 2678
      4020 ,    // 2679
      4022 ,    // 2680
      4023 ,    // 2681
      4024 ,    // 2682
      4026 ,    // 2683
      4027 ,    // 2684
      4028 ,    // 2685
      4030 ,    // 2686
      4031 ,    // 2687
      4032 ,    // 2688
      4034 ,    // 2689
      4035 ,    // 2690
      4037 ,    // 2691
      4038 ,    // 2692
      4039 ,    // 2693
      4041 ,    // 2694
      4042 ,    // 2695
      4043 ,    // 2696
      4045 ,    // 2697
      4046 ,    // 2698
      4047 ,    // 2699
      4049 ,    // 2700
      4050 ,    // 2701
      4052 ,    // 2702
      4053 ,    // 2703
      4054 ,    // 2704
      4056 ,    // 2705
      4057 ,    // 2706
      4058 ,    // 2707
      4060 ,    // 2708
      4061 ,    // 2709
      4062 ,    // 2710
      4064 ,    // 2711
      4065 ,    // 2712
      4067 ,    // 2713
      4068 ,    // 2714
      4069 ,    // 2715
      4071 ,    // 2716
      4072 ,    // 2717
      4073 ,    // 2718
      4075 ,    // 2719
      4076 ,    // 2720
      4077 ,    // 2721
      4079 ,    // 2722
      4080 ,    // 2723
      4081 ,    // 2724
      4083 ,    // 2725
      4084 ,    // 2726
      4086 ,    // 2727
      4087 ,    // 2728
      4088 ,    // 2729
      4090 ,    // 2730
      4091 ,    // 2731
      4092 ,    // 2732
      4094 ,    // 2733
      4095 ,    // 2734
      4096 ,    // 2735
      4098 ,    // 2736
      4099 ,    // 2737
      4100 ,    // 2738
      4102 ,    // 2739
      4103 ,    // 2740
      4105 ,    // 2741
      4106 ,    // 2742
      4107 ,    // 2743
      4109 ,    // 2744
      4110 ,    // 2745
      4111 ,    // 2746
      4113 ,    // 2747
      4114 ,    // 2748
      4115 ,    // 2749
      4117 ,    // 2750
      4118 ,    // 2751
      4119 ,    // 2752
      4121 ,    // 2753
      4122 ,    // 2754
      4124 ,    // 2755
      4125 ,    // 2756
      4126 ,    // 2757
      4128 ,    // 2758
      4129 ,    // 2759
      4130 ,    // 2760
      4132 ,    // 2761
      4133 ,    // 2762
      4134 ,    // 2763
      4136 ,    // 2764
      4137 ,    // 2765
      4138 ,    // 2766
      4140 ,    // 2767
      4141 ,    // 2768
      4142 ,    // 2769
      4144 ,    // 2770
      4145 ,    // 2771
      4147 ,    // 2772
      4148 ,    // 2773
      4149 ,    // 2774
      4151 ,    // 2775
      4152 ,    // 2776
      4153 ,    // 2777
      4155 ,    // 2778
      4156 ,    // 2779
      4157 ,    // 2780
      4159 ,    // 2781
      4160 ,    // 2782
      4161 ,    // 2783
      4163 ,    // 2784
      4164 ,    // 2785
      4165 ,    // 2786
      4167 ,    // 2787
      4168 ,    // 2788
      4170 ,    // 2789
      4171 ,    // 2790
      4172 ,    // 2791
      4174 ,    // 2792
      4175 ,    // 2793
      4176 ,    // 2794
      4178 ,    // 2795
      4179 ,    // 2796
      4180 ,    // 2797
      4182 ,    // 2798
      4183 ,    // 2799
      4184 ,    // 2800
      4186 ,    // 2801
      4187 ,    // 2802
      4188 ,    // 2803
      4190 ,    // 2804
      4191 ,    // 2805
      4192 ,    // 2806
      4194 ,    // 2807
      4195 ,    // 2808
      4196 ,    // 2809
      4198 ,    // 2810
      4199 ,    // 2811
      4201 ,    // 2812
      4202 ,    // 2813
      4203 ,    // 2814
      4205 ,    // 2815
      4206 ,    // 2816
      4207 ,    // 2817
      4209 ,    // 2818
      4210 ,    // 2819
      4211 ,    // 2820
      4213 ,    // 2821
      4214 ,    // 2822
      4215 ,    // 2823
      4217 ,    // 2824
      4218 ,    // 2825
      4219 ,    // 2826
      4221 ,    // 2827
      4222 ,    // 2828
      4223 ,    // 2829
      4225 ,    // 2830
      4226 ,    // 2831
      4227 ,    // 2832
      4229 ,    // 2833
      4230 ,    // 2834
      4231 ,    // 2835
      4233 ,    // 2836
      4234 ,    // 2837
      4235 ,    // 2838
      4237 ,    // 2839
      4238 ,    // 2840
      4239 ,    // 2841
      4241 ,    // 2842
      4242 ,    // 2843
      4244 ,    // 2844
      4245 ,    // 2845
      4246 ,    // 2846
      4248 ,    // 2847
      4249 ,    // 2848
      4250 ,    // 2849
      4252 ,    // 2850
      4253 ,    // 2851
      4254 ,    // 2852
      4256 ,    // 2853
      4257 ,    // 2854
      4258 ,    // 2855
      4260 ,    // 2856
      4261 ,    // 2857
      4262 ,    // 2858
      4264 ,    // 2859
      4265 ,    // 2860
      4266 ,    // 2861
      4268 ,    // 2862
      4269 ,    // 2863
      4270 ,    // 2864
      4272 ,    // 2865
      4273 ,    // 2866
      4274 ,    // 2867
      4276 ,    // 2868
      4277 ,    // 2869
      4278 ,    // 2870
      4280 ,    // 2871
      4281 ,    // 2872
      4282 ,    // 2873
      4284 ,    // 2874
      4285 ,    // 2875
      4286 ,    // 2876
      4288 ,    // 2877
      4289 ,    // 2878
      4290 ,    // 2879
      4292 ,    // 2880
      4293 ,    // 2881
      4294 ,    // 2882
      4296 ,    // 2883
      4297 ,    // 2884
      4298 ,    // 2885
      4300 ,    // 2886
      4301 ,    // 2887
      4302 ,    // 2888
      4304 ,    // 2889
      4305 ,    // 2890
      4306 ,    // 2891
      4308 ,    // 2892
      4309 ,    // 2893
      4310 ,    // 2894
      4312 ,    // 2895
      4313 ,    // 2896
      4314 ,    // 2897
      4316 ,    // 2898
      4317 ,    // 2899
      4318 ,    // 2900
      4320 ,    // 2901
      4321 ,    // 2902
      4322 ,    // 2903
      4324 ,    // 2904
      4325 ,    // 2905
      4326 ,    // 2906
      4328 ,    // 2907
      4329 ,    // 2908
      4330 ,    // 2909
      4332 ,    // 2910
      4333 ,    // 2911
      4334 ,    // 2912
      4336 ,    // 2913
      4337 ,    // 2914
      4338 ,    // 2915
      4340 ,    // 2916
      4341 ,    // 2917
      4342 ,    // 2918
      4344 ,    // 2919
      4345 ,    // 2920
      4346 ,    // 2921
      4348 ,    // 2922
      4349 ,    // 2923
      4350 ,    // 2924
      4352 ,    // 2925
      4353 ,    // 2926
      4354 ,    // 2927
      4356 ,    // 2928
      4357 ,    // 2929
      4358 ,    // 2930
      4360 ,    // 2931
      4361 ,    // 2932
      4362 ,    // 2933
      4364 ,    // 2934
      4365 ,    // 2935
      4366 ,    // 2936
      4368 ,    // 2937
      4369 ,    // 2938
      4370 ,    // 2939
      4372 ,    // 2940
      4373 ,    // 2941
      4374 ,    // 2942
      4376 ,    // 2943
      4377 ,    // 2944
      4378 ,    // 2945
      4379 ,    // 2946
      4381 ,    // 2947
      4382 ,    // 2948
      4383 ,    // 2949
      4385 ,    // 2950
      4386 ,    // 2951
      4387 ,    // 2952
      4389 ,    // 2953
      4390 ,    // 2954
      4391 ,    // 2955
      4393 ,    // 2956
      4394 ,    // 2957
      4395 ,    // 2958
      4397 ,    // 2959
      4398 ,    // 2960
      4399 ,    // 2961
      4401 ,    // 2962
      4402 ,    // 2963
      4403 ,    // 2964
      4405 ,    // 2965
      4406 ,    // 2966
      4407 ,    // 2967
      4409 ,    // 2968
      4410 ,    // 2969
      4411 ,    // 2970
      4413 ,    // 2971
      4414 ,    // 2972
      4415 ,    // 2973
      4417 ,    // 2974
      4418 ,    // 2975
      4419 ,    // 2976
      4420 ,    // 2977
      4422 ,    // 2978
      4423 ,    // 2979
      4424 ,    // 2980
      4426 ,    // 2981
      4427 ,    // 2982
      4428 ,    // 2983
      4430 ,    // 2984
      4431 ,    // 2985
      4432 ,    // 2986
      4434 ,    // 2987
      4435 ,    // 2988
      4436 ,    // 2989
      4438 ,    // 2990
      4439 ,    // 2991
      4440 ,    // 2992
      4442 ,    // 2993
      4443 ,    // 2994
      4444 ,    // 2995
      4446 ,    // 2996
      4447 ,    // 2997
      4448 ,    // 2998
      4449 ,    // 2999
      4451 ,    // 3000
      4452 ,    // 3001
      4453 ,    // 3002
      4455 ,    // 3003
      4456 ,    // 3004
      4457 ,    // 3005
      4459 ,    // 3006
      4460 ,    // 3007
      4461 ,    // 3008
      4463 ,    // 3009
      4464 ,    // 3010
      4465 ,    // 3011
      4467 ,    // 3012
      4468 ,    // 3013
      4469 ,    // 3014
      4471 ,    // 3015
      4472 ,    // 3016
      4473 ,    // 3017
      4474 ,    // 3018
      4476 ,    // 3019
      4477 ,    // 3020
      4478 ,    // 3021
      4480 ,    // 3022
      4481 ,    // 3023
      4482 ,    // 3024
      4484 ,    // 3025
      4485 ,    // 3026
      4486 ,    // 3027
      4488 ,    // 3028
      4489 ,    // 3029
      4490 ,    // 3030
      4492 ,    // 3031
      4493 ,    // 3032
      4494 ,    // 3033
      4495 ,    // 3034
      4497 ,    // 3035
      4498 ,    // 3036
      4499 ,    // 3037
      4501 ,    // 3038
      4502 ,    // 3039
      4503 ,    // 3040
      4505 ,    // 3041
      4506 ,    // 3042
      4507 ,    // 3043
      4509 ,    // 3044
      4510 ,    // 3045
      4511 ,    // 3046
      4512 ,    // 3047
      4514 ,    // 3048
      4515 ,    // 3049
      4516 ,    // 3050
      4518 ,    // 3051
      4519 ,    // 3052
      4520 ,    // 3053
      4522 ,    // 3054
      4523 ,    // 3055
      4524 ,    // 3056
      4526 ,    // 3057
      4527 ,    // 3058
      4528 ,    // 3059
      4529 ,    // 3060
      4531 ,    // 3061
      4532 ,    // 3062
      4533 ,    // 3063
      4535 ,    // 3064
      4536 ,    // 3065
      4537 ,    // 3066
      4539 ,    // 3067
      4540 ,    // 3068
      4541 ,    // 3069
      4543 ,    // 3070
      4544 ,    // 3071
      4545 ,    // 3072
      4546 ,    // 3073
      4548 ,    // 3074
      4549 ,    // 3075
      4550 ,    // 3076
      4552 ,    // 3077
      4553 ,    // 3078
      4554 ,    // 3079
      4556 ,    // 3080
      4557 ,    // 3081
      4558 ,    // 3082
      4559 ,    // 3083
      4561 ,    // 3084
      4562 ,    // 3085
      4563 ,    // 3086
      4565 ,    // 3087
      4566 ,    // 3088
      4567 ,    // 3089
      4569 ,    // 3090
      4570 ,    // 3091
      4571 ,    // 3092
      4573 ,    // 3093
      4574 ,    // 3094
      4575 ,    // 3095
      4576 ,    // 3096
      4578 ,    // 3097
      4579 ,    // 3098
      4580 ,    // 3099
      4582 ,    // 3100
      4583 ,    // 3101
      4584 ,    // 3102
      4586 ,    // 3103
      4587 ,    // 3104
      4588 ,    // 3105
      4589 ,    // 3106
      4591 ,    // 3107
      4592 ,    // 3108
      4593 ,    // 3109
      4595 ,    // 3110
      4596 ,    // 3111
      4597 ,    // 3112
      4598 ,    // 3113
      4600 ,    // 3114
      4601 ,    // 3115
      4602 ,    // 3116
      4604 ,    // 3117
      4605 ,    // 3118
      4606 ,    // 3119
      4608 ,    // 3120
      4609 ,    // 3121
      4610 ,    // 3122
      4611 ,    // 3123
      4613 ,    // 3124
      4614 ,    // 3125
      4615 ,    // 3126
      4617 ,    // 3127
      4618 ,    // 3128
      4619 ,    // 3129
      4621 ,    // 3130
      4622 ,    // 3131
      4623 ,    // 3132
      4624 ,    // 3133
      4626 ,    // 3134
      4627 ,    // 3135
      4628 ,    // 3136
      4630 ,    // 3137
      4631 ,    // 3138
      4632 ,    // 3139
      4633 ,    // 3140
      4635 ,    // 3141
      4636 ,    // 3142
      4637 ,    // 3143
      4639 ,    // 3144
      4640 ,    // 3145
      4641 ,    // 3146
      4643 ,    // 3147
      4644 ,    // 3148
      4645 ,    // 3149
      4646 ,    // 3150
      4648 ,    // 3151
      4649 ,    // 3152
      4650 ,    // 3153
      4652 ,    // 3154
      4653 ,    // 3155
      4654 ,    // 3156
      4655 ,    // 3157
      4657 ,    // 3158
      4658 ,    // 3159
      4659 ,    // 3160
      4661 ,    // 3161
      4662 ,    // 3162
      4663 ,    // 3163
      4664 ,    // 3164
      4666 ,    // 3165
      4667 ,    // 3166
      4668 ,    // 3167
      4670 ,    // 3168
      4671 ,    // 3169
      4672 ,    // 3170
      4673 ,    // 3171
      4675 ,    // 3172
      4676 ,    // 3173
      4677 ,    // 3174
      4679 ,    // 3175
      4680 ,    // 3176
      4681 ,    // 3177
      4682 ,    // 3178
      4684 ,    // 3179
      4685 ,    // 3180
      4686 ,    // 3181
      4688 ,    // 3182
      4689 ,    // 3183
      4690 ,    // 3184
      4691 ,    // 3185
      4693 ,    // 3186
      4694 ,    // 3187
      4695 ,    // 3188
      4697 ,    // 3189
      4698 ,    // 3190
      4699 ,    // 3191
      4700 ,    // 3192
      4702 ,    // 3193
      4703 ,    // 3194
      4704 ,    // 3195
      4706 ,    // 3196
      4707 ,    // 3197
      4708 ,    // 3198
      4709 ,    // 3199
      4711 ,    // 3200
      4712 ,    // 3201
      4713 ,    // 3202
      4715 ,    // 3203
      4716 ,    // 3204
      4717 ,    // 3205
      4718 ,    // 3206
      4720 ,    // 3207
      4721 ,    // 3208
      4722 ,    // 3209
      4724 ,    // 3210
      4725 ,    // 3211
      4726 ,    // 3212
      4727 ,    // 3213
      4729 ,    // 3214
      4730 ,    // 3215
      4731 ,    // 3216
      4733 ,    // 3217
      4734 ,    // 3218
      4735 ,    // 3219
      4736 ,    // 3220
      4738 ,    // 3221
      4739 ,    // 3222
      4740 ,    // 3223
      4741 ,    // 3224
      4743 ,    // 3225
      4744 ,    // 3226
      4745 ,    // 3227
      4747 ,    // 3228
      4748 ,    // 3229
      4749 ,    // 3230
      4750 ,    // 3231
      4752 ,    // 3232
      4753 ,    // 3233
      4754 ,    // 3234
      4756 ,    // 3235
      4757 ,    // 3236
      4758 ,    // 3237
      4759 ,    // 3238
      4761 ,    // 3239
      4762 ,    // 3240
      4763 ,    // 3241
      4764 ,    // 3242
      4766 ,    // 3243
      4767 ,    // 3244
      4768 ,    // 3245
      4770 ,    // 3246
      4771 ,    // 3247
      4772 ,    // 3248
      4773 ,    // 3249
      4775 ,    // 3250
      4776 ,    // 3251
      4777 ,    // 3252
      4778 ,    // 3253
      4780 ,    // 3254
      4781 ,    // 3255
      4782 ,    // 3256
      4784 ,    // 3257
      4785 ,    // 3258
      4786 ,    // 3259
      4787 ,    // 3260
      4789 ,    // 3261
      4790 ,    // 3262
      4791 ,    // 3263
      4792 ,    // 3264
      4794 ,    // 3265
      4795 ,    // 3266
      4796 ,    // 3267
      4798 ,    // 3268
      4799 ,    // 3269
      4800 ,    // 3270
      4801 ,    // 3271
      4803 ,    // 3272
      4804 ,    // 3273
      4805 ,    // 3274
      4806 ,    // 3275
      4808 ,    // 3276
      4809 ,    // 3277
      4810 ,    // 3278
      4811 ,    // 3279
      4813 ,    // 3280
      4814 ,    // 3281
      4815 ,    // 3282
      4817 ,    // 3283
      4818 ,    // 3284
      4819 ,    // 3285
      4820 ,    // 3286
      4822 ,    // 3287
      4823 ,    // 3288
      4824 ,    // 3289
      4825 ,    // 3290
      4827 ,    // 3291
      4828 ,    // 3292
      4829 ,    // 3293
      4831 ,    // 3294
      4832 ,    // 3295
      4833 ,    // 3296
      4834 ,    // 3297
      4836 ,    // 3298
      4837 ,    // 3299
      4838 ,    // 3300
      4839 ,    // 3301
      4841 ,    // 3302
      4842 ,    // 3303
      4843 ,    // 3304
      4844 ,    // 3305
      4846 ,    // 3306
      4847 ,    // 3307
      4848 ,    // 3308
      4849 ,    // 3309
      4851 ,    // 3310
      4852 ,    // 3311
      4853 ,    // 3312
      4855 ,    // 3313
      4856 ,    // 3314
      4857 ,    // 3315
      4858 ,    // 3316
      4860 ,    // 3317
      4861 ,    // 3318
      4862 ,    // 3319
      4863 ,    // 3320
      4865 ,    // 3321
      4866 ,    // 3322
      4867 ,    // 3323
      4868 ,    // 3324
      4870 ,    // 3325
      4871 ,    // 3326
      4872 ,    // 3327
      4873 ,    // 3328
      4875 ,    // 3329
      4876 ,    // 3330
      4877 ,    // 3331
      4878 ,    // 3332
      4880 ,    // 3333
      4881 ,    // 3334
      4882 ,    // 3335
      4884 ,    // 3336
      4885 ,    // 3337
      4886 ,    // 3338
      4887 ,    // 3339
      4889 ,    // 3340
      4890 ,    // 3341
      4891 ,    // 3342
      4892 ,    // 3343
      4894 ,    // 3344
      4895 ,    // 3345
      4896 ,    // 3346
      4897 ,    // 3347
      4899 ,    // 3348
      4900 ,    // 3349
      4901 ,    // 3350
      4902 ,    // 3351
      4904 ,    // 3352
      4905 ,    // 3353
      4906 ,    // 3354
      4907 ,    // 3355
      4909 ,    // 3356
      4910 ,    // 3357
      4911 ,    // 3358
      4912 ,    // 3359
      4914 ,    // 3360
      4915 ,    // 3361
      4916 ,    // 3362
      4917 ,    // 3363
      4919 ,    // 3364
      4920 ,    // 3365
      4921 ,    // 3366
      4922 ,    // 3367
      4924 ,    // 3368
      4925 ,    // 3369
      4926 ,    // 3370
      4927 ,    // 3371
      4929 ,    // 3372
      4930 ,    // 3373
      4931 ,    // 3374
      4932 ,    // 3375
      4934 ,    // 3376
      4935 ,    // 3377
      4936 ,    // 3378
      4937 ,    // 3379
      4939 ,    // 3380
      4940 ,    // 3381
      4941 ,    // 3382
      4942 ,    // 3383
      4944 ,    // 3384
      4945 ,    // 3385
      4946 ,    // 3386
      4947 ,    // 3387
      4949 ,    // 3388
      4950 ,    // 3389
      4951 ,    // 3390
      4952 ,    // 3391
      4954 ,    // 3392
      4955 ,    // 3393
      4956 ,    // 3394
      4957 ,    // 3395
      4959 ,    // 3396
      4960 ,    // 3397
      4961 ,    // 3398
      4962 ,    // 3399
      4964 ,    // 3400
      4965 ,    // 3401
      4966 ,    // 3402
      4967 ,    // 3403
      4969 ,    // 3404
      4970 ,    // 3405
      4971 ,    // 3406
      4972 ,    // 3407
      4974 ,    // 3408
      4975 ,    // 3409
      4976 ,    // 3410
      4977 ,    // 3411
      4979 ,    // 3412
      4980 ,    // 3413
      4981 ,    // 3414
      4982 ,    // 3415
      4984 ,    // 3416
      4985 ,    // 3417
      4986 ,    // 3418
      4987 ,    // 3419
      4989 ,    // 3420
      4990 ,    // 3421
      4991 ,    // 3422
      4992 ,    // 3423
      4994 ,    // 3424
      4995 ,    // 3425
      4996 ,    // 3426
      4997 ,    // 3427
      4999 ,    // 3428
      5000 ,    // 3429
      5001 ,    // 3430
      5002 ,    // 3431
      5004 ,    // 3432
      5005 ,    // 3433
      5006 ,    // 3434
      5007 ,    // 3435
      5008 ,    // 3436
      5010 ,    // 3437
      5011 ,    // 3438
      5012 ,    // 3439
      5013 ,    // 3440
      5015 ,    // 3441
      5016 ,    // 3442
      5017 ,    // 3443
      5018 ,    // 3444
      5020 ,    // 3445
      5021 ,    // 3446
      5022 ,    // 3447
      5023 ,    // 3448
      5025 ,    // 3449
      5026 ,    // 3450
      5027 ,    // 3451
      5028 ,    // 3452
      5030 ,    // 3453
      5031 ,    // 3454
      5032 ,    // 3455
      5033 ,    // 3456
      5034 ,    // 3457
      5036 ,    // 3458
      5037 ,    // 3459
      5038 ,    // 3460
      5039 ,    // 3461
      5041 ,    // 3462
      5042 ,    // 3463
      5043 ,    // 3464
      5044 ,    // 3465
      5046 ,    // 3466
      5047 ,    // 3467
      5048 ,    // 3468
      5049 ,    // 3469
      5051 ,    // 3470
      5052 ,    // 3471
      5053 ,    // 3472
      5054 ,    // 3473
      5055 ,    // 3474
      5057 ,    // 3475
      5058 ,    // 3476
      5059 ,    // 3477
      5060 ,    // 3478
      5062 ,    // 3479
      5063 ,    // 3480
      5064 ,    // 3481
      5065 ,    // 3482
      5067 ,    // 3483
      5068 ,    // 3484
      5069 ,    // 3485
      5070 ,    // 3486
      5071 ,    // 3487
      5073 ,    // 3488
      5074 ,    // 3489
      5075 ,    // 3490
      5076 ,    // 3491
      5078 ,    // 3492
      5079 ,    // 3493
      5080 ,    // 3494
      5081 ,    // 3495
      5083 ,    // 3496
      5084 ,    // 3497
      5085 ,    // 3498
      5086 ,    // 3499
      5087 ,    // 3500
      5089 ,    // 3501
      5090 ,    // 3502
      5091 ,    // 3503
      5092 ,    // 3504
      5094 ,    // 3505
      5095 ,    // 3506
      5096 ,    // 3507
      5097 ,    // 3508
      5099 ,    // 3509
      5100 ,    // 3510
      5101 ,    // 3511
      5102 ,    // 3512
      5103 ,    // 3513
      5105 ,    // 3514
      5106 ,    // 3515
      5107 ,    // 3516
      5108 ,    // 3517
      5110 ,    // 3518
      5111 ,    // 3519
      5112 ,    // 3520
      5113 ,    // 3521
      5114 ,    // 3522
      5116 ,    // 3523
      5117 ,    // 3524
      5118 ,    // 3525
      5119 ,    // 3526
      5121 ,    // 3527
      5122 ,    // 3528
      5123 ,    // 3529
      5124 ,    // 3530
      5125 ,    // 3531
      5127 ,    // 3532
      5128 ,    // 3533
      5129 ,    // 3534
      5130 ,    // 3535
      5132 ,    // 3536
      5133 ,    // 3537
      5134 ,    // 3538
      5135 ,    // 3539
      5136 ,    // 3540
      5138 ,    // 3541
      5139 ,    // 3542
      5140 ,    // 3543
      5141 ,    // 3544
      5143 ,    // 3545
      5144 ,    // 3546
      5145 ,    // 3547
      5146 ,    // 3548
      5147 ,    // 3549
      5149 ,    // 3550
      5150 ,    // 3551
      5151 ,    // 3552
      5152 ,    // 3553
      5154 ,    // 3554
      5155 ,    // 3555
      5156 ,    // 3556
      5157 ,    // 3557
      5158 ,    // 3558
      5160 ,    // 3559
      5161 ,    // 3560
      5162 ,    // 3561
      5163 ,    // 3562
      5165 ,    // 3563
      5166 ,    // 3564
      5167 ,    // 3565
      5168 ,    // 3566
      5169 ,    // 3567
      5171 ,    // 3568
      5172 ,    // 3569
      5173 ,    // 3570
      5174 ,    // 3571
      5175 ,    // 3572
      5177 ,    // 3573
      5178 ,    // 3574
      5179 ,    // 3575
      5180 ,    // 3576
      5182 ,    // 3577
      5183 ,    // 3578
      5184 ,    // 3579
      5185 ,    // 3580
      5186 ,    // 3581
      5188 ,    // 3582
      5189 ,    // 3583
      5190 ,    // 3584
      5191 ,    // 3585
      5192 ,    // 3586
      5194 ,    // 3587
      5195 ,    // 3588
      5196 ,    // 3589
      5197 ,    // 3590
      5198 ,    // 3591
      5200 ,    // 3592
      5201 ,    // 3593
      5202 ,    // 3594
      5203 ,    // 3595
      5205 ,    // 3596
      5206 ,    // 3597
      5207 ,    // 3598
      5208 ,    // 3599
      5209 ,    // 3600
      5211 ,    // 3601
      5212 ,    // 3602
      5213 ,    // 3603
      5214 ,    // 3604
      5215 ,    // 3605
      5217 ,    // 3606
      5218 ,    // 3607
      5219 ,    // 3608
      5220 ,    // 3609
      5221 ,    // 3610
      5223 ,    // 3611
      5224 ,    // 3612
      5225 ,    // 3613
      5226 ,    // 3614
      5228 ,    // 3615
      5229 ,    // 3616
      5230 ,    // 3617
      5231 ,    // 3618
      5232 ,    // 3619
      5234 ,    // 3620
      5235 ,    // 3621
      5236 ,    // 3622
      5237 ,    // 3623
      5238 ,    // 3624
      5240 ,    // 3625
      5241 ,    // 3626
      5242 ,    // 3627
      5243 ,    // 3628
      5244 ,    // 3629
      5246 ,    // 3630
      5247 ,    // 3631
      5248 ,    // 3632
      5249 ,    // 3633
      5250 ,    // 3634
      5252 ,    // 3635
      5253 ,    // 3636
      5254 ,    // 3637
      5255 ,    // 3638
      5256 ,    // 3639
      5258 ,    // 3640
      5259 ,    // 3641
      5260 ,    // 3642
      5261 ,    // 3643
      5262 ,    // 3644
      5264 ,    // 3645
      5265 ,    // 3646
      5266 ,    // 3647
      5267 ,    // 3648
      5268 ,    // 3649
      5270 ,    // 3650
      5271 ,    // 3651
      5272 ,    // 3652
      5273 ,    // 3653
      5274 ,    // 3654
      5276 ,    // 3655
      5277 ,    // 3656
      5278 ,    // 3657
      5279 ,    // 3658
      5280 ,    // 3659
      5282 ,    // 3660
      5283 ,    // 3661
      5284 ,    // 3662
      5285 ,    // 3663
      5286 ,    // 3664
      5288 ,    // 3665
      5289 ,    // 3666
      5290 ,    // 3667
      5291 ,    // 3668
      5292 ,    // 3669
      5294 ,    // 3670
      5295 ,    // 3671
      5296 ,    // 3672
      5297 ,    // 3673
      5298 ,    // 3674
      5300 ,    // 3675
      5301 ,    // 3676
      5302 ,    // 3677
      5303 ,    // 3678
      5304 ,    // 3679
      5306 ,    // 3680
      5307 ,    // 3681
      5308 ,    // 3682
      5309 ,    // 3683
      5310 ,    // 3684
      5312 ,    // 3685
      5313 ,    // 3686
      5314 ,    // 3687
      5315 ,    // 3688
      5316 ,    // 3689
      5317 ,    // 3690
      5319 ,    // 3691
      5320 ,    // 3692
      5321 ,    // 3693
      5322 ,    // 3694
      5323 ,    // 3695
      5325 ,    // 3696
      5326 ,    // 3697
      5327 ,    // 3698
      5328 ,    // 3699
      5329 ,    // 3700
      5331 ,    // 3701
      5332 ,    // 3702
      5333 ,    // 3703
      5334 ,    // 3704
      5335 ,    // 3705
      5337 ,    // 3706
      5338 ,    // 3707
      5339 ,    // 3708
      5340 ,    // 3709
      5341 ,    // 3710
      5342 ,    // 3711
      5344 ,    // 3712
      5345 ,    // 3713
      5346 ,    // 3714
      5347 ,    // 3715
      5348 ,    // 3716
      5350 ,    // 3717
      5351 ,    // 3718
      5352 ,    // 3719
      5353 ,    // 3720
      5354 ,    // 3721
      5356 ,    // 3722
      5357 ,    // 3723
      5358 ,    // 3724
      5359 ,    // 3725
      5360 ,    // 3726
      5361 ,    // 3727
      5363 ,    // 3728
      5364 ,    // 3729
      5365 ,    // 3730
      5366 ,    // 3731
      5367 ,    // 3732
      5369 ,    // 3733
      5370 ,    // 3734
      5371 ,    // 3735
      5372 ,    // 3736
      5373 ,    // 3737
      5374 ,    // 3738
      5376 ,    // 3739
      5377 ,    // 3740
      5378 ,    // 3741
      5379 ,    // 3742
      5380 ,    // 3743
      5382 ,    // 3744
      5383 ,    // 3745
      5384 ,    // 3746
      5385 ,    // 3747
      5386 ,    // 3748
      5387 ,    // 3749
      5389 ,    // 3750
      5390 ,    // 3751
      5391 ,    // 3752
      5392 ,    // 3753
      5393 ,    // 3754
      5395 ,    // 3755
      5396 ,    // 3756
      5397 ,    // 3757
      5398 ,    // 3758
      5399 ,    // 3759
      5400 ,    // 3760
      5402 ,    // 3761
      5403 ,    // 3762
      5404 ,    // 3763
      5405 ,    // 3764
      5406 ,    // 3765
      5408 ,    // 3766
      5409 ,    // 3767
      5410 ,    // 3768
      5411 ,    // 3769
      5412 ,    // 3770
      5413 ,    // 3771
      5415 ,    // 3772
      5416 ,    // 3773
      5417 ,    // 3774
      5418 ,    // 3775
      5419 ,    // 3776
      5420 ,    // 3777
      5422 ,    // 3778
      5423 ,    // 3779
      5424 ,    // 3780
      5425 ,    // 3781
      5426 ,    // 3782
      5427 ,    // 3783
      5429 ,    // 3784
      5430 ,    // 3785
      5431 ,    // 3786
      5432 ,    // 3787
      5433 ,    // 3788
      5435 ,    // 3789
      5436 ,    // 3790
      5437 ,    // 3791
      5438 ,    // 3792
      5439 ,    // 3793
      5440 ,    // 3794
      5442 ,    // 3795
      5443 ,    // 3796
      5444 ,    // 3797
      5445 ,    // 3798
      5446 ,    // 3799
      5447 ,    // 3800
      5449 ,    // 3801
      5450 ,    // 3802
      5451 ,    // 3803
      5452 ,    // 3804
      5453 ,    // 3805
      5454 ,    // 3806
      5456 ,    // 3807
      5457 ,    // 3808
      5458 ,    // 3809
      5459 ,    // 3810
      5460 ,    // 3811
      5461 ,    // 3812
      5463 ,    // 3813
      5464 ,    // 3814
      5465 ,    // 3815
      5466 ,    // 3816
      5467 ,    // 3817
      5468 ,    // 3818
      5470 ,    // 3819
      5471 ,    // 3820
      5472 ,    // 3821
      5473 ,    // 3822
      5474 ,    // 3823
      5475 ,    // 3824
      5477 ,    // 3825
      5478 ,    // 3826
      5479 ,    // 3827
      5480 ,    // 3828
      5481 ,    // 3829
      5482 ,    // 3830
      5484 ,    // 3831
      5485 ,    // 3832
      5486 ,    // 3833
      5487 ,    // 3834
      5488 ,    // 3835
      5489 ,    // 3836
      5491 ,    // 3837
      5492 ,    // 3838
      5493 ,    // 3839
      5494 ,    // 3840
      5495 ,    // 3841
      5496 ,    // 3842
      5498 ,    // 3843
      5499 ,    // 3844
      5500 ,    // 3845
      5501 ,    // 3846
      5502 ,    // 3847
      5503 ,    // 3848
      5505 ,    // 3849
      5506 ,    // 3850
      5507 ,    // 3851
      5508 ,    // 3852
      5509 ,    // 3853
      5510 ,    // 3854
      5511 ,    // 3855
      5513 ,    // 3856
      5514 ,    // 3857
      5515 ,    // 3858
      5516 ,    // 3859
      5517 ,    // 3860
      5518 ,    // 3861
      5520 ,    // 3862
      5521 ,    // 3863
      5522 ,    // 3864
      5523 ,    // 3865
      5524 ,    // 3866
      5525 ,    // 3867
      5527 ,    // 3868
      5528 ,    // 3869
      5529 ,    // 3870
      5530 ,    // 3871
      5531 ,    // 3872
      5532 ,    // 3873
      5533 ,    // 3874
      5535 ,    // 3875
      5536 ,    // 3876
      5537 ,    // 3877
      5538 ,    // 3878
      5539 ,    // 3879
      5540 ,    // 3880
      5542 ,    // 3881
      5543 ,    // 3882
      5544 ,    // 3883
      5545 ,    // 3884
      5546 ,    // 3885
      5547 ,    // 3886
      5548 ,    // 3887
      5550 ,    // 3888
      5551 ,    // 3889
      5552 ,    // 3890
      5553 ,    // 3891
      5554 ,    // 3892
      5555 ,    // 3893
      5557 ,    // 3894

      5558 ,    // 3895
      5559 ,    // 3896
      5560 ,    // 3897
      5561 ,    // 3898
      5562 ,    // 3899
      5563 ,    // 3900
      5565 ,    // 3901
      5566 ,    // 3902
      5567 ,    // 3903
      5568 ,    // 3904
      5569 ,    // 3905
      5570 ,    // 3906
      5571 ,    // 3907
      5573 ,    // 3908
      5574 ,    // 3909
      5575 ,    // 3910
      5576 ,    // 3911
      5577 ,    // 3912
      5578 ,    // 3913
      5580 ,    // 3914
      5581 ,    // 3915
      5582 ,    // 3916
      5583 ,    // 3917
      5584 ,    // 3918
      5585 ,    // 3919
      5586 ,    // 3920
      5588 ,    // 3921
      5589 ,    // 3922
      5590 ,    // 3923
      5591 ,    // 3924
      5592 ,    // 3925
      5593 ,    // 3926
      5594 ,    // 3927
      5596 ,    // 3928
      5597 ,    // 3929
      5598 ,    // 3930
      5599 ,    // 3931
      5600 ,    // 3932
      5601 ,    // 3933
      5602 ,    // 3934
      5604 ,    // 3935
      5605 ,    // 3936
      5606 ,    // 3937
      5607 ,    // 3938
      5608 ,    // 3939
      5609 ,    // 3940
      5610 ,    // 3941
      5612 ,    // 3942
      5613 ,    // 3943
      5614 ,    // 3944
      5615 ,    // 3945
      5616 ,    // 3946
      5617 ,    // 3947
      5618 ,    // 3948
      5620 ,    // 3949
      5621 ,    // 3950
      5622 ,    // 3951
      5623 ,    // 3952
      5624 ,    // 3953
      5625 ,    // 3954
      5626 ,    // 3955
      5628 ,    // 3956
      5629 ,    // 3957
      5630 ,    // 3958
      5631 ,    // 3959
      5632 ,    // 3960
      5633 ,    // 3961
      5634 ,    // 3962
      5635 ,    // 3963
      5637 ,    // 3964
      5638 ,    // 3965
      5639 ,    // 3966
      5640 ,    // 3967
      5641 ,    // 3968
      5642 ,    // 3969
      5643 ,    // 3970
      5645 ,    // 3971
      5646 ,    // 3972
      5647 ,    // 3973
      5648 ,    // 3974
      5649 ,    // 3975
      5650 ,    // 3976
      5651 ,    // 3977
      5653 ,    // 3978
      5654 ,    // 3979
      5655 ,    // 3980
      5656 ,    // 3981
      5657 ,    // 3982
      5658 ,    // 3983
      5659 ,    // 3984
      5660 ,    // 3985
      5662 ,    // 3986
      5663 ,    // 3987
      5664 ,    // 3988
      5665 ,    // 3989
      5666 ,    // 3990
      5667 ,    // 3991
      5668 ,    // 3992
      5670 ,    // 3993
      5671 ,    // 3994
      5672 ,    // 3995
      5673 ,    // 3996
      5674 ,    // 3997
      5675 ,    // 3998
      5676 ,    // 3999
      5677 ,    // 4000
      5679 ,    // 4001
      5680 ,    // 4002
      5681 ,    // 4003
      5682 ,    // 4004
      5683 ,    // 4005
      5684 ,    // 4006
      5685 ,    // 4007
      5686 ,    // 4008
      5688 ,    // 4009
      5689 ,    // 4010
      5690 ,    // 4011
      5691 ,    // 4012
      5692 ,    // 4013
      5693 ,    // 4014
      5694 ,    // 4015
      5695 ,    // 4016
      5697 ,    // 4017
      5698 ,    // 4018
      5699 ,    // 4019
      5700 ,    // 4020
      5701 ,    // 4021
      5702 ,    // 4022
      5703 ,    // 4023
      5704 ,    // 4024
      5706 ,    // 4025
      5707 ,    // 4026
      5708 ,    // 4027
      5709 ,    // 4028
      5710 ,    // 4029
      5711 ,    // 4030
      5712 ,    // 4031
      5713 ,    // 4032
      5715 ,    // 4033
      5716 ,    // 4034
      5717 ,    // 4035
      5718 ,    // 4036
      5719 ,    // 4037
      5720 ,    // 4038
      5721 ,    // 4039
      5722 ,    // 4040
      5724 ,    // 4041
      5725 ,    // 4042
      5726 ,    // 4043
      5727 ,    // 4044
      5728 ,    // 4045
      5729 ,    // 4046
      5730 ,    // 4047
      5731 ,    // 4048
      5733 ,    // 4049
      5734 ,    // 4050
      5735 ,    // 4051
      5736 ,    // 4052
      5737 ,    // 4053
      5738 ,    // 4054
      5739 ,    // 4055
      5740 ,    // 4056
      5741 ,    // 4057
      5743 ,    // 4058
      5744 ,    // 4059
      5745 ,    // 4060
      5746 ,    // 4061
      5747 ,    // 4062
      5748 ,    // 4063
      5749 ,    // 4064
      5750 ,    // 4065
      5752 ,    // 4066
      5753 ,    // 4067
      5754 ,    // 4068
      5755 ,    // 4069
      5756 ,    // 4070
      5757 ,    // 4071
      5758 ,    // 4072
      5759 ,    // 4073
      5760 ,    // 4074
      5762 ,    // 4075
      5763 ,    // 4076
      5764 ,    // 4077
      5765 ,    // 4078
      5766 ,    // 4079
      5767 ,    // 4080
      5768 ,    // 4081
      5769 ,    // 4082
      5770 ,    // 4083
      5772 ,    // 4084
      5773 ,    // 4085
      5774 ,    // 4086
      5775 ,    // 4087
      5776 ,    // 4088
      5777 ,    // 4089
      5778 ,    // 4090
      5779 ,    // 4091
      5780 ,    // 4092
      5782 ,    // 4093
      5783 ,    // 4094
      5784 ,    // 4095
      5785 ,    // 4096
      5786 ,    // 4097
      5787 ,    // 4098
      5788 ,    // 4099
      5789 ,    // 4100
      5790 ,    // 4101
      5792 ,    // 4102
      5793 ,    // 4103
      5794 ,    // 4104
      5795 ,    // 4105
      5796 ,    // 4106
      5797 ,    // 4107
      5798 ,    // 4108
      5799 ,    // 4109
      5800 ,    // 4110
      5801 ,    // 4111
      5803 ,    // 4112
      5804 ,    // 4113
      5805 ,    // 4114
      5806 ,    // 4115
      5807 ,    // 4116
      5808 ,    // 4117
      5809 ,    // 4118
      5810 ,    // 4119
      5811 ,    // 4120
      5813 ,    // 4121
      5814 ,    // 4122
      5815 ,    // 4123
      5816 ,    // 4124
      5817 ,    // 4125
      5818 ,    // 4126
      5819 ,    // 4127
      5820 ,    // 4128
      5821 ,    // 4129
      5822 ,    // 4130
      5824 ,    // 4131
      5825 ,    // 4132
      5826 ,    // 4133
      5827 ,    // 4134
      5828 ,    // 4135
      5829 ,    // 4136
      5830 ,    // 4137
      5831 ,    // 4138
      5832 ,    // 4139
      5833 ,    // 4140
      5835 ,    // 4141
      5836 ,    // 4142
      5837 ,    // 4143
      5838 ,    // 4144
      5839 ,    // 4145
      5840 ,    // 4146
      5841 ,    // 4147
      5842 ,    // 4148
      5843 ,    // 4149
      5844 ,    // 4150
      5846 ,    // 4151
      5847 ,    // 4152
      5848 ,    // 4153
      5849 ,    // 4154
      5850 ,    // 4155
      5851 ,    // 4156
      5852 ,    // 4157
      5853 ,    // 4158
      5854 ,    // 4159
      5855 ,    // 4160
      5857 ,    // 4161
      5858 ,    // 4162
      5859 ,    // 4163
      5860 ,    // 4164
      5861 ,    // 4165
      5862 ,    // 4166
      5863 ,    // 4167
      5864 ,    // 4168
      5865 ,    // 4169
      5866 ,    // 4170
      5867 ,    // 4171
      5869 ,    // 4172
      5870 ,    // 4173
      5871 ,    // 4174
      5872 ,    // 4175
      5873 ,    // 4176
      5874 ,    // 4177
      5875 ,    // 4178
      5876 ,    // 4179
      5877 ,    // 4180
      5878 ,    // 4181
      5879 ,    // 4182
      5881 ,    // 4183
      5882 ,    // 4184
      5883 ,    // 4185
      5884 ,    // 4186
      5885 ,    // 4187
      5886 ,    // 4188
      5887 ,    // 4189
      5888 ,    // 4190
      5889 ,    // 4191
      5890 ,    // 4192
      5891 ,    // 4193
      5893 ,    // 4194
      5894 ,    // 4195
      5895 ,    // 4196
      5896 ,    // 4197
      5897 ,    // 4198
      5898 ,    // 4199
      5899 ,    // 4200
      5900 ,    // 4201
      5901 ,    // 4202
      5902 ,    // 4203
      5903 ,    // 4204
      5905 ,    // 4205
      5906 ,    // 4206
      5907 ,    // 4207
      5908 ,    // 4208
      5909 ,    // 4209
      5910 ,    // 4210
      5911 ,    // 4211
      5912 ,    // 4212
      5913 ,    // 4213
      5914 ,    // 4214
      5915 ,    // 4215
      5916 ,    // 4216
      5918 ,    // 4217
      5919 ,    // 4218
      5920 ,    // 4219
      5921 ,    // 4220
      5922 ,    // 4221
      5923 ,    // 4222
      5924 ,    // 4223
      5925 ,    // 4224
      5926 ,    // 4225
      5927 ,    // 4226
      5928 ,    // 4227
      5929 ,    // 4228
      5931 ,    // 4229
      5932 ,    // 4230
      5933 ,    // 4231
      5934 ,    // 4232
      5935 ,    // 4233
      5936 ,    // 4234
      5937 ,    // 4235
      5938 ,    // 4236
      5939 ,    // 4237
      5940 ,    // 4238
      5941 ,    // 4239
      5942 ,    // 4240
      5943 ,    // 4241
      5945 ,    // 4242
      5946 ,    // 4243
      5947 ,    // 4244
      5948 ,    // 4245
      5949 ,    // 4246
      5950 ,    // 4247
      5951 ,    // 4248
      5952 ,    // 4249
      5953 ,    // 4250
      5954 ,    // 4251
      5955 ,    // 4252
      5956 ,    // 4253
      5957 ,    // 4254
      5959 ,    // 4255
      5960 ,    // 4256
      5961 ,    // 4257
      5962 ,    // 4258
      5963 ,    // 4259
      5964 ,    // 4260
      5965 ,    // 4261
      5966 ,    // 4262
      5967 ,    // 4263
      5968 ,    // 4264
      5969 ,    // 4265
      5970 ,    // 4266
      5971 ,    // 4267
      5972 ,    // 4268
      5974 ,    // 4269
      5975 ,    // 4270
      5976 ,    // 4271
      5977 ,    // 4272
      5978 ,    // 4273
      5979 ,    // 4274
      5980 ,    // 4275
      5981 ,    // 4276
      5982 ,    // 4277
      5983 ,    // 4278
      5984 ,    // 4279
      5985 ,    // 4280
      5986 ,    // 4281
      5987 ,    // 4282
      5989 ,    // 4283
      5990 ,    // 4284
      5991 ,    // 4285
      5992 ,    // 4286
      5993 ,    // 4287
      5994 ,    // 4288
      5995 ,    // 4289
      5996 ,    // 4290
      5997 ,    // 4291
      5998 ,    // 4292
      5999 ,    // 4293
      6000 ,    // 4294
      6001 ,    // 4295
      6002 ,    // 4296
      6003 ,    // 4297
      6005 ,    // 4298
      6006 ,    // 4299
      6007 ,    // 4300
      6008 ,    // 4301
      6009 ,    // 4302
      6010 ,    // 4303
      6011 ,    // 4304
      6012 ,    // 4305
      6013 ,    // 4306
      6014 ,    // 4307
      6015 ,    // 4308
      6016 ,    // 4309
      6017 ,    // 4310
      6018 ,    // 4311
      6019 ,    // 4312
      6021 ,    // 4313
      6022 ,    // 4314
      6023 ,    // 4315
      6024 ,    // 4316
      6025 ,    // 4317
      6026 ,    // 4318
      6027 ,    // 4319
      6028 ,    // 4320
      6029 ,    // 4321
      6030 ,    // 4322
      6031 ,    // 4323
      6032 ,    // 4324
      6033 ,    // 4325
      6034 ,    // 4326
      6035 ,    // 4327
      6036 ,    // 4328
      6037 ,    // 4329
      6039 ,    // 4330
      6040 ,    // 4331
      6041 ,    // 4332
      6042 ,    // 4333
      6043 ,    // 4334
      6044 ,    // 4335
      6045 ,    // 4336
      6046 ,    // 4337
      6047 ,    // 4338
      6048 ,    // 4339
      6049 ,    // 4340
      6050 ,    // 4341
      6051 ,    // 4342
      6052 ,    // 4343
      6053 ,    // 4344
      6054 ,    // 4345
      6055 ,    // 4346
      6056 ,    // 4347
      6058 ,    // 4348
      6059 ,    // 4349
      6060 ,    // 4350
      6061 ,    // 4351
      6062 ,    // 4352
      6063 ,    // 4353
      6064 ,    // 4354
      6065 ,    // 4355
      6066 ,    // 4356
      6067 ,    // 4357
      6068 ,    // 4358
      6069 ,    // 4359
      6070 ,    // 4360
      6071 ,    // 4361
      6072 ,    // 4362
      6073 ,    // 4363
      6074 ,    // 4364
      6075 ,    // 4365
      6076 ,    // 4366
      6078 ,    // 4367
      6079 ,    // 4368
      6080 ,    // 4369
      6081 ,    // 4370
      6082 ,    // 4371
      6083 ,    // 4372
      6084 ,    // 4373
      6085 ,    // 4374
      6086 ,    // 4375
      6087 ,    // 4376
      6088 ,    // 4377
      6089 ,    // 4378
      6090 ,    // 4379
      6091 ,    // 4380
      6092 ,    // 4381
      6093 ,    // 4382
      6094 ,    // 4383
      6095 ,    // 4384
      6096 ,    // 4385
      6097 ,    // 4386
      6099 ,    // 4387
      6100 ,    // 4388
      6101 ,    // 4389
      6102 ,    // 4390
      6103 ,    // 4391
      6104 ,    // 4392
      6105 ,    // 4393
      6106 ,    // 4394
      6107 ,    // 4395
      6108 ,    // 4396
      6109 ,    // 4397
      6110 ,    // 4398
      6111 ,    // 4399
      6112 ,    // 4400
      6113 ,    // 4401
      6114 ,    // 4402
      6115 ,    // 4403
      6116 ,    // 4404
      6117 ,    // 4405
      6118 ,    // 4406
      6119 ,    // 4407
      6120 ,    // 4408
      6121 ,    // 4409
      6122 ,    // 4410
      6124 ,    // 4411
      6125 ,    // 4412
      6126 ,    // 4413
      6127 ,    // 4414
      6128 ,    // 4415
      6129 ,    // 4416
      6130 ,    // 4417
      6131 ,    // 4418
      6132 ,    // 4419
      6133 ,    // 4420
      6134 ,    // 4421
      6135 ,    // 4422
      6136 ,    // 4423
      6137 ,    // 4424
      6138 ,    // 4425
      6139 ,    // 4426
      6140 ,    // 4427
      6141 ,    // 4428
      6142 ,    // 4429
      6143 ,    // 4430
      6144 ,    // 4431
      6145 ,    // 4432
      6146 ,    // 4433
      6147 ,    // 4434
      6148 ,    // 4435
      6149 ,    // 4436
      6151 ,    // 4437
      6152 ,    // 4438
      6153 ,    // 4439
      6154 ,    // 4440
      6155 ,    // 4441
      6156 ,    // 4442
      6157 ,    // 4443
      6158 ,    // 4444
      6159 ,    // 4445
      6160 ,    // 4446
      6161 ,    // 4447
      6162 ,    // 4448
      6163 ,    // 4449
      6164 ,    // 4450
      6165 ,    // 4451
      6166 ,    // 4452
      6167 ,    // 4453
      6168 ,    // 4454
      6169 ,    // 4455
      6170 ,    // 4456
      6171 ,    // 4457
      6172 ,    // 4458
      6173 ,    // 4459
      6174 ,    // 4460
      6175 ,    // 4461
      6176 ,    // 4462
      6177 ,    // 4463
      6178 ,    // 4464
      6179 ,    // 4465
      6180 ,    // 4466
      6181 ,    // 4467
      6182 ,    // 4468
      6183 ,    // 4469
      6185 ,    // 4470
      6186 ,    // 4471
      6187 ,    // 4472
      6188 ,    // 4473
      6189 ,    // 4474
      6190 ,    // 4475
      6191 ,    // 4476
      6192 ,    // 4477
      6193 ,    // 4478
      6194 ,    // 4479
      6195 ,    // 4480
      6196 ,    // 4481
      6197 ,    // 4482
      6198 ,    // 4483
      6199 ,    // 4484
      6200 ,    // 4485
      6201 ,    // 4486
      6202 ,    // 4487
      6203 ,    // 4488
      6204 ,    // 4489
      6205 ,    // 4490
      6206 ,    // 4491
      6207 ,    // 4492
      6208 ,    // 4493
      6209 ,    // 4494
      6210 ,    // 4495
      6211 ,    // 4496
      6212 ,    // 4497
      6213 ,    // 4498
      6214 ,    // 4499
      6215 ,    // 4500
      6216 ,    // 4501
      6217 ,    // 4502
      6218 ,    // 4503
      6219 ,    // 4504
      6220 ,    // 4505
      6221 ,    // 4506
      6222 ,    // 4507
      6223 ,    // 4508
      6224 ,    // 4509
      6225 ,    // 4510
      6226 ,    // 4511
      6227 ,    // 4512
      6228 ,    // 4513
      6229 ,    // 4514
      6230 ,    // 4515
      6232 ,    // 4516
      6233 ,    // 4517
      6234 ,    // 4518
      6235 ,    // 4519
      6236 ,    // 4520
      6237 ,    // 4521
      6238 ,    // 4522
      6239 ,    // 4523
      6240 ,    // 4524
      6241 ,    // 4525
      6242 ,    // 4526
      6243 ,    // 4527
      6244 ,    // 4528
      6245 ,    // 4529
      6246 ,    // 4530
      6247 ,    // 4531
      6248 ,    // 4532
      6249 ,    // 4533
      6250 ,    // 4534
      6251 ,    // 4535
      6252 ,    // 4536
      6253 ,    // 4537
      6254 ,    // 4538
      6255 ,    // 4539
      6256 ,    // 4540
      6257 ,    // 4541
      6258 ,    // 4542
      6259 ,    // 4543
      6260 ,    // 4544
      6261 ,    // 4545
      6262 ,    // 4546
      6263 ,    // 4547
      6264 ,    // 4548
      6265 ,    // 4549
      6266 ,    // 4550
      6267 ,    // 4551
      6268 ,    // 4552
      6269 ,    // 4553
      6270 ,    // 4554
      6271 ,    // 4555
      6272 ,    // 4556
      6273 ,    // 4557
      6274 ,    // 4558
      6275 ,    // 4559
      6276 ,    // 4560
      6277 ,    // 4561
      6278 ,    // 4562
      6279 ,    // 4563
      6280 ,    // 4564
      6281 ,    // 4565
      6282 ,    // 4566
      6283 ,    // 4567
      6284 ,    // 4568
      6285 ,    // 4569
      6286 ,    // 4570
      6287 ,    // 4571
      6288 ,    // 4572
      6289 ,    // 4573
      6290 ,    // 4574
      6291 ,    // 4575
      6292 ,    // 4576
      6293 ,    // 4577
      6294 ,    // 4578
      6295 ,    // 4579
      6296 ,    // 4580
      6297 ,    // 4581
      6298 ,    // 4582
      6299 ,    // 4583
      6300 ,    // 4584
      6301 ,    // 4585
      6302 ,    // 4586
      6303 ,    // 4587
      6304 ,    // 4588
      6305 ,    // 4589
      6306 ,    // 4590
      6307 ,    // 4591
      6308 ,    // 4592
      6309 ,    // 4593
      6310 ,    // 4594
      6311 ,    // 4595
      6312 ,    // 4596
      6313 ,    // 4597
      6314 ,    // 4598
      6315 ,    // 4599
      6316 ,    // 4600
      6317 ,    // 4601
      6318 ,    // 4602
      6319 ,    // 4603
      6320 ,    // 4604
      6321 ,    // 4605
      6322 ,    // 4606
      6323 ,    // 4607
      6324 ,    // 4608
      6325 ,    // 4609
      6326 ,    // 4610
      6327 ,    // 4611
      6328 ,    // 4612
      6329 ,    // 4613
      6330 ,    // 4614
      6331 ,    // 4615
      6332 ,    // 4616
      6333 ,    // 4617
      6334 ,    // 4618
      6335 ,    // 4619
      6336 ,    // 4620
      6337 ,    // 4621
      6338 ,    // 4622
      6339 ,    // 4623
      6340 ,    // 4624
      6341 ,    // 4625
      6342 ,    // 4626
      6343 ,    // 4627
      6344 ,    // 4628
      6345 ,    // 4629
      6346 ,    // 4630
      6347 ,    // 4631
      6348 ,    // 4632
      6349 ,    // 4633
      6350 ,    // 4634
      6351 ,    // 4635
      6352 ,    // 4636
      6353 ,    // 4637
      6354 ,    // 4638
      6355 ,    // 4639
      6356 ,    // 4640
      6357 ,    // 4641
      6358 ,    // 4642
      6359 ,    // 4643
      6360 ,    // 4644
      6361 ,    // 4645
      6362 ,    // 4646
      6363 ,    // 4647
      6364 ,    // 4648
      6365 ,    // 4649
      6366 ,    // 4650
      6367 ,    // 4651
      6368 ,    // 4652
      6369 ,    // 4653
      6370 ,    // 4654
      6371 ,    // 4655
      6372 ,    // 4656
      6373 ,    // 4657
      6374 ,    // 4658
      6374 ,    // 4659
      6375 ,    // 4660
      6376 ,    // 4661
      6377 ,    // 4662
      6378 ,    // 4663
      6379 ,    // 4664
      6380 ,    // 4665
      6381 ,    // 4666
      6382 ,    // 4667
      6383 ,    // 4668
      6384 ,    // 4669
      6385 ,    // 4670
      6386 ,    // 4671
      6387 ,    // 4672
      6388 ,    // 4673
      6389 ,    // 4674
      6390 ,    // 4675
      6391 ,    // 4676
      6392 ,    // 4677
      6393 ,    // 4678
      6394 ,    // 4679
      6395 ,    // 4680
      6396 ,    // 4681
      6397 ,    // 4682
      6398 ,    // 4683
      6399 ,    // 4684
      6400 ,    // 4685
      6401 ,    // 4686
      6402 ,    // 4687
      6403 ,    // 4688
      6404 ,    // 4689
      6405 ,    // 4690
      6406 ,    // 4691
      6407 ,    // 4692
      6408 ,    // 4693
      6409 ,    // 4694
      6410 ,    // 4695
      6411 ,    // 4696
      6412 ,    // 4697
      6413 ,    // 4698
      6414 ,    // 4699
      6415 ,    // 4700
      6416 ,    // 4701
      6417 ,    // 4702
      6418 ,    // 4703
      6419 ,    // 4704
      6419 ,    // 4705
      6420 ,    // 4706
      6421 ,    // 4707
      6422 ,    // 4708
      6423 ,    // 4709
      6424 ,    // 4710
      6425 ,    // 4711
      6426 ,    // 4712
      6427 ,    // 4713
      6428 ,    // 4714
      6429 ,    // 4715
      6430 ,    // 4716
      6431 ,    // 4717
      6432 ,    // 4718
      6433 ,    // 4719
      6434 ,    // 4720
      6435 ,    // 4721
      6436 ,    // 4722
      6437 ,    // 4723
      6438 ,    // 4724
      6439 ,    // 4725
      6440 ,    // 4726
      6441 ,    // 4727
      6442 ,    // 4728
      6443 ,    // 4729
      6444 ,    // 4730
      6445 ,    // 4731
      6446 ,    // 4732
      6447 ,    // 4733
      6448 ,    // 4734
      6449 ,    // 4735
      6450 ,    // 4736
      6450 ,    // 4737
      6451 ,    // 4738
      6452 ,    // 4739
      6453 ,    // 4740
      6454 ,    // 4741
      6455 ,    // 4742
      6456 ,    // 4743
      6457 ,    // 4744
      6458 ,    // 4745
      6459 ,    // 4746
      6460 ,    // 4747
      6461 ,    // 4748
      6462 ,    // 4749
      6463 ,    // 4750
      6464 ,    // 4751
      6465 ,    // 4752
      6466 ,    // 4753
      6467 ,    // 4754
      6468 ,    // 4755
      6469 ,    // 4756
      6470 ,    // 4757
      6471 ,    // 4758
      6472 ,    // 4759
      6473 ,    // 4760
      6474 ,    // 4761
      6475 ,    // 4762
      6475 ,    // 4763
      6476 ,    // 4764
      6477 ,    // 4765
      6478 ,    // 4766
      6479 ,    // 4767
      6480 ,    // 4768
      6481 ,    // 4769
      6482 ,    // 4770
      6483 ,    // 4771
      6484 ,    // 4772
      6485 ,    // 4773
      6486 ,    // 4774
      6487 ,    // 4775
      6488 ,    // 4776
      6489 ,    // 4777
      6490 ,    // 4778
      6491 ,    // 4779
      6492 ,    // 4780
      6493 ,    // 4781
      6494 ,    // 4782
      6495 ,    // 4783
      6496 ,    // 4784
      6497 ,    // 4785
      6497 ,    // 4786
      6498 ,    // 4787
      6499 ,    // 4788
      6500 ,    // 4789
      6501 ,    // 4790
      6502 ,    // 4791
      6503 ,    // 4792
      6504 ,    // 4793
      6505 ,    // 4794
      6506 ,    // 4795
      6507 ,    // 4796
      6508 ,    // 4797
      6509 ,    // 4798
      6510 ,    // 4799
      6511 ,    // 4800
      6512 ,    // 4801
      6513 ,    // 4802
      6514 ,    // 4803
      6515 ,    // 4804
      6516 ,    // 4805
      6516 ,    // 4806
      6517 ,    // 4807
      6518 ,    // 4808
      6519 ,    // 4809
      6520 ,    // 4810
      6521 ,    // 4811
      6522 ,    // 4812
      6523 ,    // 4813
      6524 ,    // 4814
      6525 ,    // 4815
      6526 ,    // 4816
      6527 ,    // 4817
      6528 ,    // 4818
      6529 ,    // 4819
      6530 ,    // 4820
      6531 ,    // 4821
      6532 ,    // 4822
      6533 ,    // 4823
      6534 ,    // 4824
      6534 ,    // 4825
      6535 ,    // 4826
      6536 ,    // 4827
      6537 ,    // 4828
      6538 ,    // 4829
      6539 ,    // 4830
      6540 ,    // 4831
      6541 ,    // 4832
      6542 ,    // 4833
      6543 ,    // 4834
      6544 ,    // 4835
      6545 ,    // 4836
      6546 ,    // 4837
      6547 ,    // 4838
      6548 ,    // 4839
      6549 ,    // 4840
      6550 ,    // 4841
      6550 ,    // 4842
      6551 ,    // 4843
      6552 ,    // 4844
      6553 ,    // 4845
      6554 ,    // 4846
      6555 ,    // 4847
      6556 ,    // 4848
      6557 ,    // 4849
      6558 ,    // 4850
      6559 ,    // 4851
      6560 ,    // 4852
      6561 ,    // 4853
      6562 ,    // 4854
      6563 ,    // 4855
      6564 ,    // 4856
      6565 ,    // 4857
      6565 ,    // 4858
      6566 ,    // 4859
      6567 ,    // 4860
      6568 ,    // 4861
      6569 ,    // 4862
      6570 ,    // 4863
      6571 ,    // 4864
      6572 ,    // 4865
      6573 ,    // 4866
      6574 ,    // 4867
      6575 ,    // 4868
      6576 ,    // 4869
      6577 ,    // 4870
      6578 ,    // 4871
      6579 ,    // 4872
      6579 ,    // 4873
      6580 ,    // 4874
      6581 ,    // 4875
      6582 ,    // 4876
      6583 ,    // 4877
      6584 ,    // 4878
      6585 ,    // 4879
      6586 ,    // 4880
      6587 ,    // 4881
      6588 ,    // 4882
      6589 ,    // 4883
      6590 ,    // 4884
      6591 ,    // 4885
      6592 ,    // 4886
      6593 ,    // 4887
      6593 ,    // 4888
      6594 ,    // 4889
      6595 ,    // 4890
      6596 ,    // 4891
      6597 ,    // 4892
      6598 ,    // 4893
      6599 ,    // 4894
      6600 ,    // 4895
      6601 ,    // 4896
      6602 ,    // 4897
      6603 ,    // 4898
      6604 ,    // 4899
      6605 ,    // 4900
      6606 ,    // 4901
      6606 ,    // 4902
      6607 ,    // 4903
      6608 ,    // 4904
      6609 ,    // 4905
      6610 ,    // 4906
      6611 ,    // 4907
      6612 ,    // 4908
      6613 ,    // 4909
      6614 ,    // 4910
      6615 ,    // 4911
      6616 ,    // 4912
      6617 ,    // 4913
      6618 ,    // 4914
      6618 ,    // 4915
      6619 ,    // 4916
      6620 ,    // 4917
      6621 ,    // 4918
      6622 ,    // 4919
      6623 ,    // 4920
      6624 ,    // 4921
      6625 ,    // 4922
      6626 ,    // 4923
      6627 ,    // 4924
      6628 ,    // 4925
      6629 ,    // 4926
      6629 ,    // 4927
      6630 ,    // 4928
      6631 ,    // 4929
      6632 ,    // 4930
      6633 ,    // 4931
      6634 ,    // 4932
      6635 ,    // 4933
      6636 ,    // 4934
      6637 ,    // 4935
      6638 ,    // 4936
      6639 ,    // 4937
      6640 ,    // 4938
      6640 ,    // 4939
      6641 ,    // 4940
      6642 ,    // 4941
      6643 ,    // 4942
      6644 ,    // 4943
      6645 ,    // 4944
      6646 ,    // 4945
      6647 ,    // 4946
      6648 ,    // 4947
      6649 ,    // 4948
      6650 ,    // 4949
      6651 ,    // 4950
      6651 ,    // 4951
      6652 ,    // 4952
      6653 ,    // 4953
      6654 ,    // 4954
      6655 ,    // 4955
      6656 ,    // 4956
      6657 ,    // 4957
      6658 ,    // 4958
      6659 ,    // 4959
      6660 ,    // 4960
      6661 ,    // 4961
      6662 ,    // 4962
      6662 ,    // 4963
      6663 ,    // 4964
      6664 ,    // 4965
      6665 ,    // 4966
      6666 ,    // 4967
      6667 ,    // 4968
      6668 ,    // 4969
      6669 ,    // 4970
      6670 ,    // 4971
      6671 ,    // 4972
      6672 ,    // 4973
      6672 ,    // 4974
      6673 ,    // 4975
      6674 ,    // 4976
      6675 ,    // 4977
      6676 ,    // 4978
      6677 ,    // 4979
      6678 ,    // 4980
      6679 ,    // 4981
      6680 ,    // 4982
      6681 ,    // 4983
      6681 ,    // 4984
      6682 ,    // 4985
      6683 ,    // 4986
      6684 ,    // 4987
      6685 ,    // 4988
      6686 ,    // 4989
      6687 ,    // 4990
      6688 ,    // 4991
      6689 ,    // 4992
      6690 ,    // 4993
      6691 ,    // 4994
      6691 ,    // 4995
      6692 ,    // 4996
      6693 ,    // 4997
      6694 ,    // 4998
      6695 ,    // 4999
      6696 ,    // 5000
      6697 ,    // 5001
      6698 ,    // 5002
      6699 ,    // 5003
      6700 ,    // 5004
      6700 ,    // 5005
      6701 ,    // 5006
      6702 ,    // 5007
      6703 ,    // 5008
      6704 ,    // 5009
      6705 ,    // 5010
      6706 ,    // 5011
      6707 ,    // 5012
      6708 ,    // 5013
      6709 ,    // 5014
      6709 ,    // 5015
      6710 ,    // 5016
      6711 ,    // 5017
      6712 ,    // 5018
      6713 ,    // 5019
      6714 ,    // 5020
      6715 ,    // 5021
      6716 ,    // 5022
      6717 ,    // 5023
      6717 ,    // 5024
      6718 ,    // 5025
      6719 ,    // 5026
      6720 ,    // 5027
      6721 ,    // 5028
      6722 ,    // 5029
      6723 ,    // 5030
      6724 ,    // 5031
      6725 ,    // 5032
      6726 ,    // 5033
      6726 ,    // 5034
      6727 ,    // 5035
      6728 ,    // 5036
      6729 ,    // 5037
      6730 ,    // 5038
      6731 ,    // 5039
      6732 ,    // 5040
      6733 ,    // 5041
      6734 ,    // 5042
      6734 ,    // 5043
      6735 ,    // 5044
      6736 ,    // 5045
      6737 ,    // 5046
      6738 ,    // 5047
      6739 ,    // 5048
      6740 ,    // 5049
      6741 ,    // 5050
      6742 ,    // 5051
      6742 ,    // 5052
      6743 ,    // 5053
      6744 ,    // 5054
      6745 ,    // 5055
      6746 ,    // 5056
      6747 ,    // 5057
      6748 ,    // 5058
      6749 ,    // 5059
      6750 ,    // 5060
      6750 ,    // 5061
      6751 ,    // 5062
      6752 ,    // 5063
      6753 ,    // 5064
      6754 ,    // 5065
      6755 ,    // 5066
      6756 ,    // 5067
      6757 ,    // 5068
      6758 ,    // 5069
      6758 ,    // 5070
      6759 ,    // 5071
      6760 ,    // 5072
      6761 ,    // 5073
      6762 ,    // 5074
      6763 ,    // 5075
      6764 ,    // 5076
      6765 ,    // 5077
      6765 ,    // 5078
      6766 ,    // 5079
      6767 ,    // 5080
      6768 ,    // 5081
      6769 ,    // 5082
      6770 ,    // 5083
      6771 ,    // 5084
      6772 ,    // 5085
      6773 ,    // 5086
      6773 ,    // 5087
      6774 ,    // 5088
      6775 ,    // 5089
      6776 ,    // 5090
      6777 ,    // 5091
      6778 ,    // 5092
      6779 ,    // 5093
      6780 ,    // 5094
      6780 ,    // 5095
      6781 ,    // 5096
      6782 ,    // 5097
      6783 ,    // 5098
      6784 ,    // 5099
      6785 ,    // 5100
      6786 ,    // 5101
      6787 ,    // 5102
      6787 ,    // 5103
      6788 ,    // 5104
      6789 ,    // 5105
      6790 ,    // 5106
      6791 ,    // 5107
      6792 ,    // 5108
      6793 ,    // 5109
      6794 ,    // 5110
      6794 ,    // 5111
      6795 ,    // 5112
      6796 ,    // 5113
      6797 ,    // 5114
      6798 ,    // 5115
      6799 ,    // 5116
      6800 ,    // 5117
      6801 ,    // 5118
      6801 ,    // 5119
      6802 ,    // 5120
      6803 ,    // 5121
      6804 ,    // 5122
      6805 ,    // 5123
      6806 ,    // 5124
      6807 ,    // 5125
      6808 ,    // 5126
      6808 ,    // 5127
      6809 ,    // 5128
      6810 ,    // 5129
      6811 ,    // 5130
      6812 ,    // 5131
      6813 ,    // 5132
      6814 ,    // 5133
      6814 ,    // 5134
      6815 ,    // 5135
      6816 ,    // 5136
      6817 ,    // 5137
      6818 ,    // 5138
      6819 ,    // 5139
      6820 ,    // 5140
      6821 ,    // 5141
      6821 ,    // 5142
      6822 ,    // 5143
      6823 ,    // 5144
      6824 ,    // 5145
      6825 ,    // 5146
      6826 ,    // 5147
      6827 ,    // 5148
      6827 ,    // 5149
      6828 ,    // 5150
      6829 ,    // 5151
      6830 ,    // 5152
      6831 ,    // 5153
      6832 ,    // 5154
      6833 ,    // 5155
      6834 ,    // 5156
      6834 ,    // 5157
      6835 ,    // 5158
      6836 ,    // 5159
      6837 ,    // 5160
      6838 ,    // 5161
      6839 ,    // 5162
      6840 ,    // 5163
      6840 ,    // 5164
      6841 ,    // 5165
      6842 ,    // 5166
      6843 ,    // 5167
      6844 ,    // 5168
      6845 ,    // 5169
      6846 ,    // 5170
      6846 ,    // 5171
      6847 ,    // 5172
      6848 ,    // 5173
      6849 ,    // 5174
      6850 ,    // 5175
      6851 ,    // 5176
      6852 ,    // 5177
      6852 ,    // 5178
      6853 ,    // 5179
      6854 ,    // 5180
      6855 ,    // 5181
      6856 ,    // 5182
      6857 ,    // 5183
      6858 ,    // 5184
      6858 ,    // 5185
      6859 ,    // 5186
      6860 ,    // 5187
      6861 ,    // 5188
      6862 ,    // 5189
      6863 ,    // 5190
      6864 ,    // 5191
      6864 ,    // 5192
      6865 ,    // 5193
      6866 ,    // 5194
      6867 ,    // 5195
      6868 ,    // 5196
      6869 ,    // 5197
      6870 ,    // 5198
      6870 ,    // 5199
      6871 ,    // 5200
      6872 ,    // 5201
      6873 ,    // 5202
      6874 ,    // 5203
      6875 ,    // 5204
      6875 ,    // 5205
      6876 ,    // 5206
      6877 ,    // 5207
      6878 ,    // 5208
      6879 ,    // 5209
      6880 ,    // 5210
      6881 ,    // 5211
      6881 ,    // 5212
      6882 ,    // 5213
      6883 ,    // 5214
      6884 ,    // 5215
      6885 ,    // 5216
      6886 ,    // 5217
      6887 ,    // 5218
      6887 ,    // 5219
      6888 ,    // 5220
      6889 ,    // 5221
      6890 ,    // 5222
      6891 ,    // 5223
      6892 ,    // 5224
      6892 ,    // 5225
      6893 ,    // 5226
      6894 ,    // 5227
      6895 ,    // 5228
      6896 ,    // 5229
      6897 ,    // 5230
      6897 ,    // 5231
      6898 ,    // 5232
      6899 ,    // 5233
      6900 ,    // 5234
      6901 ,    // 5235
      6902 ,    // 5236
      6903 ,    // 5237
      6903 ,    // 5238
      6904 ,    // 5239
      6905 ,    // 5240
      6906 ,    // 5241
      6907 ,    // 5242
      6908 ,    // 5243
      6908 ,    // 5244
      6909 ,    // 5245
      6910 ,    // 5246
      6911 ,    // 5247
      6912 ,    // 5248
      6913 ,    // 5249
      6913 ,    // 5250
      6914 ,    // 5251
      6915 ,    // 5252
      6916 ,    // 5253
      6917 ,    // 5254
      6918 ,    // 5255
      6919 ,    // 5256
      6919 ,    // 5257
      6920 ,    // 5258
      6921 ,    // 5259
      6922 ,    // 5260
      6923 ,    // 5261
      6924 ,    // 5262
      6924 ,    // 5263
      6925 ,    // 5264
      6926 ,    // 5265
      6927 ,    // 5266
      6928 ,    // 5267
      6929 ,    // 5268
      6929 ,    // 5269
      6930 ,    // 5270
      6931 ,    // 5271
      6932 ,    // 5272
      6933 ,    // 5273
      6934 ,    // 5274
      6934 ,    // 5275
      6935 ,    // 5276
      6936 ,    // 5277
      6937 ,    // 5278
      6938 ,    // 5279
      6939 ,    // 5280
      6939 ,    // 5281
      6940 ,    // 5282
      6941 ,    // 5283
      6942 ,    // 5284
      6943 ,    // 5285
      6944 ,    // 5286
      6944 ,    // 5287
      6945 ,    // 5288
      6946 ,    // 5289
      6947 ,    // 5290
      6948 ,    // 5291
      6948 ,    // 5292
      6949 ,    // 5293
      6950 ,    // 5294
      6951 ,    // 5295
      6952 ,    // 5296
      6953 ,    // 5297
      6953 ,    // 5298
      6954 ,    // 5299
      6955 ,    // 5300
      6956 ,    // 5301
      6957 ,    // 5302
      6958 ,    // 5303
      6958 ,    // 5304
      6959 ,    // 5305
      6960 ,    // 5306
      6961 ,    // 5307
      6962 ,    // 5308
      6963 ,    // 5309
      6963 ,    // 5310
      6964 ,    // 5311
      6965 ,    // 5312
      6966 ,    // 5313
      6967 ,    // 5314
      6967 ,    // 5315
      6968 ,    // 5316
      6969 ,    // 5317
      6970 ,    // 5318
      6971 ,    // 5319
      6972 ,    // 5320
      6972 ,    // 5321
      6973 ,    // 5322
      6974 ,    // 5323
      6975 ,    // 5324
      6976 ,    // 5325
      6976 ,    // 5326
      6977 ,    // 5327
      6978 ,    // 5328
      6979 ,    // 5329
      6980 ,    // 5330
      6981 ,    // 5331
      6981 ,    // 5332
      6982 ,    // 5333
      6983 ,    // 5334
      6984 ,    // 5335
      6985 ,    // 5336
      6985 ,    // 5337
      6986 ,    // 5338
      6987 ,    // 5339
      6988 ,    // 5340
      6989 ,    // 5341
      6990 ,    // 5342
      6990 ,    // 5343
      6991 ,    // 5344
      6992 ,    // 5345
      6993 ,    // 5346
      6994 ,    // 5347
      6994 ,    // 5348
      6995 ,    // 5349
      6996 ,    // 5350
      6997 ,    // 5351
      6998 ,    // 5352
      6999 ,    // 5353
      6999 ,    // 5354
      7000 ,    // 5355
      7001 ,    // 5356
      7002 ,    // 5357
      7003 ,    // 5358
      7003 ,    // 5359
      7004 ,    // 5360
      7005 ,    // 5361
      7006 ,    // 5362
      7007 ,    // 5363
      7007 ,    // 5364
      7008 ,    // 5365
      7009 ,    // 5366
      7010 ,    // 5367
      7011 ,    // 5368
      7011 ,    // 5369
      7012 ,    // 5370
      7013 ,    // 5371
      7014 ,    // 5372
      7015 ,    // 5373
      7016 ,    // 5374
      7016 ,    // 5375
      7017 ,    // 5376
      7018 ,    // 5377
      7019 ,    // 5378
      7020 ,    // 5379
      7020 ,    // 5380
      7021 ,    // 5381
      7022 ,    // 5382
      7023 ,    // 5383
      7024 ,    // 5384
      7024 ,    // 5385
      7025 ,    // 5386
      7026 ,    // 5387
      7027 ,    // 5388
      7028 ,    // 5389
      7028 ,    // 5390
      7029 ,    // 5391
      7030 ,    // 5392
      7031 ,    // 5393
      7032 ,    // 5394
      7032 ,    // 5395
      7033 ,    // 5396
      7034 ,    // 5397
      7035 ,    // 5398
      7036 ,    // 5399
      7036 ,    // 5400
      7037 ,    // 5401
      7038 ,    // 5402
      7039 ,    // 5403
      7040 ,    // 5404
      7040 ,    // 5405
      7041 ,    // 5406
      7042 ,    // 5407
      7043 ,    // 5408
      7044 ,    // 5409
      7044 ,    // 5410
      7045 ,    // 5411
      7046 ,    // 5412
      7047 ,    // 5413
      7048 ,    // 5414
      7048 ,    // 5415
      7049 ,    // 5416
      7050 ,    // 5417
      7051 ,    // 5418
      7052 ,    // 5419
      7052 ,    // 5420
      7053 ,    // 5421
      7054 ,    // 5422
      7055 ,    // 5423
      7056 ,    // 5424
      7056 ,    // 5425
      7057 ,    // 5426
      7058 ,    // 5427
      7059 ,    // 5428
      7060 ,    // 5429
      7060 ,    // 5430
      7061 ,    // 5431
      7062 ,    // 5432
      7063 ,    // 5433
      7063 ,    // 5434
      7064 ,    // 5435
      7065 ,    // 5436
      7066 ,    // 5437
      7067 ,    // 5438
      7067 ,    // 5439
      7068 ,    // 5440
      7069 ,    // 5441
      7070 ,    // 5442
      7071 ,    // 5443
      7071 ,    // 5444
      7072 ,    // 5445
      7073 ,    // 5446
      7074 ,    // 5447
      7075 ,    // 5448
      7075 ,    // 5449
      7076 ,    // 5450
      7077 ,    // 5451
      7078 ,    // 5452
      7078 ,    // 5453
      7079 ,    // 5454
      7080 ,    // 5455
      7081 ,    // 5456
      7082 ,    // 5457
      7082 ,    // 5458
      7083 ,    // 5459
      7084 ,    // 5460
      7085 ,    // 5461
      7086 ,    // 5462
      7086 ,    // 5463
      7087 ,    // 5464
      7088 ,    // 5465
      7089 ,    // 5466
      7089 ,    // 5467
      7090 ,    // 5468
      7091 ,    // 5469
      7092 ,    // 5470
      7093 ,    // 5471
      7093 ,    // 5472
      7094 ,    // 5473
      7095 ,    // 5474
      7096 ,    // 5475
      7096 ,    // 5476
      7097 ,    // 5477
      7098 ,    // 5478
      7099 ,    // 5479
      7100 ,    // 5480
      7100 ,    // 5481
      7101 ,    // 5482
      7102 ,    // 5483
      7103 ,    // 5484
      7103 ,    // 5485
      7104 ,    // 5486
      7105 ,    // 5487
      7106 ,    // 5488
      7107 ,    // 5489
      7107 ,    // 5490
      7108 ,    // 5491
      7109 ,    // 5492
      7110 ,    // 5493
      7110 ,    // 5494
      7111 ,    // 5495
      7112 ,    // 5496
      7113 ,    // 5497
      7114 ,    // 5498
      7114 ,    // 5499
      7115 ,    // 5500
      7116 ,    // 5501
      7117 ,    // 5502
      7117 ,    // 5503
      7118 ,    // 5504
      7119 ,    // 5505
      7120 ,    // 5506
      7121 ,    // 5507
      7121 ,    // 5508
      7122 ,    // 5509
      7123 ,    // 5510
      7124 ,    // 5511
      7124 ,    // 5512
      7125 ,    // 5513
      7126 ,    // 5514
      7127 ,    // 5515
      7127 ,    // 5516
      7128 ,    // 5517
      7129 ,    // 5518
      7130 ,    // 5519
      7131 ,    // 5520
      7131 ,    // 5521
      7132 ,    // 5522
      7133 ,    // 5523
      7134 ,    // 5524
      7134 ,    // 5525
      7135 ,    // 5526
      7136 ,    // 5527
      7137 ,    // 5528
      7137 ,    // 5529
      7138 ,    // 5530
      7139 ,    // 5531
      7140 ,    // 5532
      7141 ,    // 5533
      7141 ,    // 5534
      7142 ,    // 5535
      7143 ,    // 5536
      7144 ,    // 5537
      7144 ,    // 5538
      7145 ,    // 5539
      7146 ,    // 5540
      7147 ,    // 5541
      7147 ,    // 5542
      7148 ,    // 5543
      7149 ,    // 5544
      7150 ,    // 5545
      7150 ,    // 5546
      7151 ,    // 5547
      7152 ,    // 5548
      7153 ,    // 5549
      7154 ,    // 5550
      7154 ,    // 5551
      7155 ,    // 5552
      7156 ,    // 5553
      7157 ,    // 5554
      7157 ,    // 5555
      7158 ,    // 5556
      7159 ,    // 5557
      7160 ,    // 5558
      7160 ,    // 5559
      7161 ,    // 5560
      7162 ,    // 5561
      7163 ,    // 5562
      7163 ,    // 5563
      7164 ,    // 5564
      7165 ,    // 5565
      7166 ,    // 5566
      7166 ,    // 5567
      7167 ,    // 5568
      7168 ,    // 5569
      7169 ,    // 5570
      7169 ,    // 5571
      7170 ,    // 5572
      7171 ,    // 5573
      7172 ,    // 5574
      7172 ,    // 5575
      7173 ,    // 5576
      7174 ,    // 5577
      7175 ,    // 5578
      7175 ,    // 5579
      7176 ,    // 5580
      7177 ,    // 5581
      7178 ,    // 5582
      7179 ,    // 5583
      7179 ,    // 5584
      7180 ,    // 5585
      7181 ,    // 5586
      7182 ,    // 5587
      7182 ,    // 5588
      7183 ,    // 5589
      7184 ,    // 5590
      7185 ,    // 5591
      7185 ,    // 5592
      7186 ,    // 5593
      7187 ,    // 5594
      7188 ,    // 5595
      7188 ,    // 5596
      7189 ,    // 5597
      7190 ,    // 5598
      7191 ,    // 5599
      7191 ,    // 5600
      7192 ,    // 5601
      7193 ,    // 5602
      7193 ,    // 5603
      7194 ,    // 5604
      7195 ,    // 5605
      7196 ,    // 5606
      7196 ,    // 5607
      7197 ,    // 5608
      7198 ,    // 5609
      7199 ,    // 5610
      7199 ,    // 5611
      7200 ,    // 5612
      7201 ,    // 5613
      7202 ,    // 5614
      7202 ,    // 5615
      7203 ,    // 5616
      7204 ,    // 5617
      7205 ,    // 5618
      7205 ,    // 5619
      7206 ,    // 5620
      7207 ,    // 5621
      7208 ,    // 5622
      7208 ,    // 5623
      7209 ,    // 5624
      7210 ,    // 5625
      7211 ,    // 5626
      7211 ,    // 5627
      7212 ,    // 5628
      7213 ,    // 5629
      7214 ,    // 5630
      7214 ,    // 5631
      7215 ,    // 5632
      7216 ,    // 5633
      7217 ,    // 5634
      7217 ,    // 5635
      7218 ,    // 5636
      7219 ,    // 5637
      7219 ,    // 5638
      7220 ,    // 5639
      7221 ,    // 5640
      7222 ,    // 5641
      7222 ,    // 5642
      7223 ,    // 5643
      7224 ,    // 5644
      7225 ,    // 5645
      7225 ,    // 5646
      7226 ,    // 5647
      7227 ,    // 5648
      7228 ,    // 5649
      7228 ,    // 5650
      7229 ,    // 5651
      7230 ,    // 5652
      7231 ,    // 5653
      7231 ,    // 5654
      7232 ,    // 5655
      7233 ,    // 5656
      7233 ,    // 5657
      7234 ,    // 5658
      7235 ,    // 5659
      7236 ,    // 5660
      7236 ,    // 5661
      7237 ,    // 5662
      7238 ,    // 5663
      7239 ,    // 5664
      7239 ,    // 5665
      7240 ,    // 5666
      7241 ,    // 5667
      7242 ,    // 5668
      7242 ,    // 5669
      7243 ,    // 5670
      7244 ,    // 5671
      7244 ,    // 5672
      7245 ,    // 5673
      7246 ,    // 5674
      7247 ,    // 5675
      7247 ,    // 5676
      7248 ,    // 5677
      7249 ,    // 5678
      7250 ,    // 5679
      7250 ,    // 5680
      7251 ,    // 5681
      7252 ,    // 5682
      7252 ,    // 5683
      7253 ,    // 5684
      7254 ,    // 5685
      7255 ,    // 5686
      7255 ,    // 5687
      7256 ,    // 5688
      7257 ,    // 5689
      7257 ,    // 5690
      7258 ,    // 5691
      7259 ,    // 5692
      7260 ,    // 5693
      7260 ,    // 5694
      7261 ,    // 5695
      7262 ,    // 5696
      7263 ,    // 5697
      7263 ,    // 5698
      7264 ,    // 5699
      7265 ,    // 5700
      7265 ,    // 5701
      7266 ,    // 5702
      7267 ,    // 5703
      7268 ,    // 5704
      7268 ,    // 5705
      7269 ,    // 5706
      7270 ,    // 5707
      7270 ,    // 5708
      7271 ,    // 5709
      7272 ,    // 5710
      7273 ,    // 5711
      7273 ,    // 5712
      7274 ,    // 5713
      7275 ,    // 5714
      7276 ,    // 5715
      7276 ,    // 5716
      7277 ,    // 5717
      7278 ,    // 5718
      7278 ,    // 5719
      7279 ,    // 5720
      7280 ,    // 5721
      7281 ,    // 5722
      7281 ,    // 5723
      7282 ,    // 5724
      7283 ,    // 5725
      7283 ,    // 5726
      7284 ,    // 5727
      7285 ,    // 5728
      7286 ,    // 5729
      7286 ,    // 5730
      7287 ,    // 5731
      7288 ,    // 5732
      7288 ,    // 5733
      7289 ,    // 5734
      7290 ,    // 5735
      7291 ,    // 5736
      7291 ,    // 5737
      7292 ,    // 5738
      7293 ,    // 5739
      7293 ,    // 5740
      7294 ,    // 5741
      7295 ,    // 5742
      7295 ,    // 5743
      7296 ,    // 5744
      7297 ,    // 5745
      7298 ,    // 5746
      7298 ,    // 5747
      7299 ,    // 5748
      7300 ,    // 5749
      7300 ,    // 5750
      7301 ,    // 5751
      7302 ,    // 5752
      7303 ,    // 5753
      7303 ,    // 5754
      7304 ,    // 5755
      7305 ,    // 5756
      7305 ,    // 5757
      7306 ,    // 5758
      7307 ,    // 5759
      7308 ,    // 5760
      7308 ,    // 5761
      7309 ,    // 5762
      7310 ,    // 5763
      7310 ,    // 5764
      7311 ,    // 5765
      7312 ,    // 5766
      7312 ,    // 5767
      7313 ,    // 5768
      7314 ,    // 5769
      7315 ,    // 5770
      7315 ,    // 5771
      7316 ,    // 5772
      7317 ,    // 5773
      7317 ,    // 5774
      7318 ,    // 5775
      7319 ,    // 5776
      7319 ,    // 5777
      7320 ,    // 5778
      7321 ,    // 5779
      7322 ,    // 5780
      7322 ,    // 5781
      7323 ,    // 5782
      7324 ,    // 5783
      7324 ,    // 5784
      7325 ,    // 5785
      7326 ,    // 5786
      7326 ,    // 5787
      7327 ,    // 5788
      7328 ,    // 5789
      7329 ,    // 5790
      7329 ,    // 5791
      7330 ,    // 5792
      7331 ,    // 5793
      7331 ,    // 5794
      7332 ,    // 5795
      7333 ,    // 5796
      7333 ,    // 5797
      7334 ,    // 5798
      7335 ,    // 5799
      7336 ,    // 5800
      7336 ,    // 5801
      7337 ,    // 5802
      7338 ,    // 5803
      7338 ,    // 5804
      7339 ,    // 5805
      7340 ,    // 5806
      7340 ,    // 5807
      7341 ,    // 5808
      7342 ,    // 5809
      7342 ,    // 5810
      7343 ,    // 5811
      7344 ,    // 5812
      7345 ,    // 5813
      7345 ,    // 5814
      7346 ,    // 5815
      7347 ,    // 5816
      7347 ,    // 5817
      7348 ,    // 5818
      7349 ,    // 5819
      7349 ,    // 5820
      7350 ,    // 5821
      7351 ,    // 5822
      7351 ,    // 5823
      7352 ,    // 5824
      7353 ,    // 5825
      7353 ,    // 5826
      7354 ,    // 5827
      7355 ,    // 5828
      7356 ,    // 5829
      7356 ,    // 5830
      7357 ,    // 5831
      7358 ,    // 5832
      7358 ,    // 5833
      7359 ,    // 5834
      7360 ,    // 5835
      7360 ,    // 5836
      7361 ,    // 5837
      7362 ,    // 5838
      7362 ,    // 5839
      7363 ,    // 5840
      7364 ,    // 5841
      7364 ,    // 5842
      7365 ,    // 5843
      7366 ,    // 5844
      7367 ,    // 5845
      7367 ,    // 5846
      7368 ,    // 5847
      7369 ,    // 5848
      7369 ,    // 5849
      7370 ,    // 5850
      7371 ,    // 5851
      7371 ,    // 5852
      7372 ,    // 5853
      7373 ,    // 5854
      7373 ,    // 5855
      7374 ,    // 5856
      7375 ,    // 5857
      7375 ,    // 5858
      7376 ,    // 5859
      7377 ,    // 5860
      7377 ,    // 5861
      7378 ,    // 5862
      7379 ,    // 5863
      7379 ,    // 5864
      7380 ,    // 5865
      7381 ,    // 5866
      7381 ,    // 5867
      7382 ,    // 5868
      7383 ,    // 5869
      7383 ,    // 5870
      7384 ,    // 5871
      7385 ,    // 5872
      7386 ,    // 5873
      7386 ,    // 5874
      7387 ,    // 5875
      7388 ,    // 5876
      7388 ,    // 5877
      7389 ,    // 5878
      7390 ,    // 5879
      7390 ,    // 5880
      7391 ,    // 5881
      7392 ,    // 5882
      7392 ,    // 5883
      7393 ,    // 5884
      7394 ,    // 5885
      7394 ,    // 5886
      7395 ,    // 5887
      7396 ,    // 5888
      7396 ,    // 5889
      7397 ,    // 5890
      7398 ,    // 5891
      7398 ,    // 5892
      7399 ,    // 5893
      7400 ,    // 5894
      7400 ,    // 5895
      7401 ,    // 5896
      7402 ,    // 5897
      7402 ,    // 5898
      7403 ,    // 5899
      7404 ,    // 5900
      7404 ,    // 5901
      7405 ,    // 5902
      7406 ,    // 5903
      7406 ,    // 5904
      7407 ,    // 5905
      7408 ,    // 5906
      7408 ,    // 5907
      7409 ,    // 5908
      7410 ,    // 5909
      7410 ,    // 5910
      7411 ,    // 5911
      7412 ,    // 5912
      7412 ,    // 5913
      7413 ,    // 5914
      7414 ,    // 5915
      7414 ,    // 5916
      7415 ,    // 5917
      7416 ,    // 5918
      7416 ,    // 5919
      7417 ,    // 5920
      7418 ,    // 5921
      7418 ,    // 5922
      7419 ,    // 5923
      7420 ,    // 5924
      7420 ,    // 5925
      7421 ,    // 5926
      7422 ,    // 5927
      7422 ,    // 5928
      7423 ,    // 5929
      7424 ,    // 5930
      7424 ,    // 5931
      7425 ,    // 5932
      7425 ,    // 5933
      7426 ,    // 5934
      7427 ,    // 5935
      7427 ,    // 5936
      7428 ,    // 5937
      7429 ,    // 5938
      7429 ,    // 5939
      7430 ,    // 5940
      7431 ,    // 5941
      7431 ,    // 5942
      7432 ,    // 5943
      7433 ,    // 5944
      7433 ,    // 5945
      7434 ,    // 5946
      7435 ,    // 5947
      7435 ,    // 5948
      7436 ,    // 5949
      7437 ,    // 5950
      7437 ,    // 5951
      7438 ,    // 5952
      7439 ,    // 5953
      7439 ,    // 5954
      7440 ,    // 5955
      7441 ,    // 5956
      7441 ,    // 5957
      7442 ,    // 5958
      7443 ,    // 5959
      7443 ,    // 5960
      7444 ,    // 5961
      7444 ,    // 5962
      7445 ,    // 5963
      7446 ,    // 5964
      7446 ,    // 5965
      7447 ,    // 5966
      7448 ,    // 5967
      7448 ,    // 5968
      7449 ,    // 5969
      7450 ,    // 5970
      7450 ,    // 5971
      7451 ,    // 5972
      7452 ,    // 5973
      7452 ,    // 5974
      7453 ,    // 5975
      7454 ,    // 5976
      7454 ,    // 5977
      7455 ,    // 5978
      7455 ,    // 5979
      7456 ,    // 5980
      7457 ,    // 5981
      7457 ,    // 5982
      7458 ,    // 5983
      7459 ,    // 5984
      7459 ,    // 5985
      7460 ,    // 5986
      7461 ,    // 5987
      7461 ,    // 5988
      7462 ,    // 5989
      7463 ,    // 5990
      7463 ,    // 5991
      7464 ,    // 5992
      7465 ,    // 5993
      7465 ,    // 5994
      7466 ,    // 5995
      7466 ,    // 5996
      7467 ,    // 5997
      7468 ,    // 5998
      7468 ,    // 5999
      7469 ,    // 6000
      7470 ,    // 6001
      7470 ,    // 6002
      7471 ,    // 6003
      7472 ,    // 6004
      7472 ,    // 6005
      7473 ,    // 6006
      7473 ,    // 6007
      7474 ,    // 6008
      7475 ,    // 6009
      7475 ,    // 6010
      7476 ,    // 6011
      7477 ,    // 6012
      7477 ,    // 6013
      7478 ,    // 6014
      7479 ,    // 6015
      7479 ,    // 6016
      7480 ,    // 6017
      7480 ,    // 6018
      7481 ,    // 6019
      7482 ,    // 6020
      7482 ,    // 6021
      7483 ,    // 6022
      7484 ,    // 6023
      7484 ,    // 6024
      7485 ,    // 6025
      7486 ,    // 6026
      7486 ,    // 6027
      7487 ,    // 6028
      7487 ,    // 6029
      7488 ,    // 6030
      7489 ,    // 6031
      7489 ,    // 6032
      7490 ,    // 6033
      7491 ,    // 6034
      7491 ,    // 6035
      7492 ,    // 6036
      7492 ,    // 6037
      7493 ,    // 6038
      7494 ,    // 6039
      7494 ,    // 6040
      7495 ,    // 6041
      7496 ,    // 6042
      7496 ,    // 6043
      7497 ,    // 6044
      7498 ,    // 6045
      7498 ,    // 6046
      7499 ,    // 6047
      7499 ,    // 6048
      7500 ,    // 6049
      7501 ,    // 6050
      7501 ,    // 6051
      7502 ,    // 6052
      7503 ,    // 6053
      7503 ,    // 6054
      7504 ,    // 6055
      7504 ,    // 6056
      7505 ,    // 6057
      7506 ,    // 6058
      7506 ,    // 6059
      7507 ,    // 6060
      7508 ,    // 6061
      7508 ,    // 6062
      7509 ,    // 6063
      7509 ,    // 6064
      7510 ,    // 6065
      7511 ,    // 6066
      7511 ,    // 6067
      7512 ,    // 6068
      7513 ,    // 6069
      7513 ,    // 6070
      7514 ,    // 6071
      7514 ,    // 6072
      7515 ,    // 6073
      7516 ,    // 6074
      7516 ,    // 6075
      7517 ,    // 6076
      7517 ,    // 6077
      7518 ,    // 6078
      7519 ,    // 6079
      7519 ,    // 6080
      7520 ,    // 6081
      7521 ,    // 6082
      7521 ,    // 6083
      7522 ,    // 6084
      7522 ,    // 6085
      7523 ,    // 6086
      7524 ,    // 6087
      7524 ,    // 6088
      7525 ,    // 6089
      7525 ,    // 6090
      7526 ,    // 6091
      7527 ,    // 6092
      7527 ,    // 6093
      7528 ,    // 6094
      7529 ,    // 6095
      7529 ,    // 6096
      7530 ,    // 6097
      7530 ,    // 6098
      7531 ,    // 6099
      7532 ,    // 6100
      7532 ,    // 6101
      7533 ,    // 6102
      7533 ,    // 6103
      7534 ,    // 6104
      7535 ,    // 6105
      7535 ,    // 6106
      7536 ,    // 6107
      7537 ,    // 6108
      7537 ,    // 6109
      7538 ,    // 6110
      7538 ,    // 6111
      7539 ,    // 6112
      7540 ,    // 6113
      7540 ,    // 6114
      7541 ,    // 6115
      7541 ,    // 6116
      7542 ,    // 6117
      7543 ,    // 6118
      7543 ,    // 6119
      7544 ,    // 6120
      7544 ,    // 6121
      7545 ,    // 6122
      7546 ,    // 6123
      7546 ,    // 6124
      7547 ,    // 6125
      7547 ,    // 6126
      7548 ,    // 6127
      7549 ,    // 6128
      7549 ,    // 6129
      7550 ,    // 6130
      7550 ,    // 6131
      7551 ,    // 6132
      7552 ,    // 6133
      7552 ,    // 6134
      7553 ,    // 6135
      7554 ,    // 6136
      7554 ,    // 6137
      7555 ,    // 6138
      7555 ,    // 6139
      7556 ,    // 6140
      7557 ,    // 6141
      7557 ,    // 6142
      7558 ,    // 6143
      7558 ,    // 6144
      7559 ,    // 6145
      7560 ,    // 6146
      7560 ,    // 6147
      7561 ,    // 6148
      7561 ,    // 6149
      7562 ,    // 6150
      7563 ,    // 6151
      7563 ,    // 6152
      7564 ,    // 6153
      7564 ,    // 6154
      7565 ,    // 6155
      7565 ,    // 6156
      7566 ,    // 6157
      7567 ,    // 6158
      7567 ,    // 6159
      7568 ,    // 6160
      7568 ,    // 6161
      7569 ,    // 6162
      7570 ,    // 6163
      7570 ,    // 6164
      7571 ,    // 6165
      7571 ,    // 6166
      7572 ,    // 6167
      7573 ,    // 6168
      7573 ,    // 6169
      7574 ,    // 6170
      7574 ,    // 6171
      7575 ,    // 6172
      7576 ,    // 6173
      7576 ,    // 6174
      7577 ,    // 6175
      7577 ,    // 6176
      7578 ,    // 6177
      7579 ,    // 6178
      7579 ,    // 6179
      7580 ,    // 6180
      7580 ,    // 6181
      7581 ,    // 6182
      7582 ,    // 6183
      7582 ,    // 6184
      7583 ,    // 6185
      7583 ,    // 6186
      7584 ,    // 6187
      7584 ,    // 6188
      7585 ,    // 6189
      7586 ,    // 6190
      7586 ,    // 6191
      7587 ,    // 6192
      7587 ,    // 6193
      7588 ,    // 6194
      7589 ,    // 6195
      7589 ,    // 6196
      7590 ,    // 6197
      7590 ,    // 6198
      7591 ,    // 6199
      7591 ,    // 6200
      7592 ,    // 6201
      7593 ,    // 6202
      7593 ,    // 6203
      7594 ,    // 6204
      7594 ,    // 6205
      7595 ,    // 6206
      7596 ,    // 6207
      7596 ,    // 6208
      7597 ,    // 6209
      7597 ,    // 6210
      7598 ,    // 6211
      7598 ,    // 6212
      7599 ,    // 6213
      7600 ,    // 6214
      7600 ,    // 6215
      7601 ,    // 6216
      7601 ,    // 6217
      7602 ,    // 6218
      7603 ,    // 6219
      7603 ,    // 6220
      7604 ,    // 6221
      7604 ,    // 6222
      7605 ,    // 6223
      7605 ,    // 6224
      7606 ,    // 6225
      7607 ,    // 6226
      7607 ,    // 6227
      7608 ,    // 6228
      7608 ,    // 6229
      7609 ,    // 6230
      7609 ,    // 6231
      7610 ,    // 6232
      7611 ,    // 6233
      7611 ,    // 6234
      7612 ,    // 6235
      7612 ,    // 6236
      7613 ,    // 6237
      7614 ,    // 6238
      7614 ,    // 6239
      7615 ,    // 6240
      7615 ,    // 6241
      7616 ,    // 6242
      7616 ,    // 6243
      7617 ,    // 6244
      7618 ,    // 6245
      7618 ,    // 6246
      7619 ,    // 6247
      7619 ,    // 6248
      7620 ,    // 6249
      7620 ,    // 6250
      7621 ,    // 6251
      7622 ,    // 6252
      7622 ,    // 6253
      7623 ,    // 6254
      7623 ,    // 6255
      7624 ,    // 6256
      7624 ,    // 6257
      7625 ,    // 6258
      7626 ,    // 6259
      7626 ,    // 6260
      7627 ,    // 6261
      7627 ,    // 6262
      7628 ,    // 6263
      7628 ,    // 6264
      7629 ,    // 6265
      7629 ,    // 6266
      7630 ,    // 6267
      7631 ,    // 6268
      7631 ,    // 6269
      7632 ,    // 6270
      7632 ,    // 6271
      7633 ,    // 6272
      7633 ,    // 6273
      7634 ,    // 6274
      7635 ,    // 6275
      7635 ,    // 6276
      7636 ,    // 6277
      7636 ,    // 6278
      7637 ,    // 6279
      7637 ,    // 6280
      7638 ,    // 6281
      7639 ,    // 6282
      7639 ,    // 6283
      7640 ,    // 6284
      7640 ,    // 6285
      7641 ,    // 6286
      7641 ,    // 6287
      7642 ,    // 6288
      7642 ,    // 6289
      7643 ,    // 6290
      7644 ,    // 6291
      7644 ,    // 6292
      7645 ,    // 6293
      7645 ,    // 6294
      7646 ,    // 6295
      7646 ,    // 6296
      7647 ,    // 6297
      7647 ,    // 6298
      7648 ,    // 6299
      7649 ,    // 6300
      7649 ,    // 6301
      7650 ,    // 6302
      7650 ,    // 6303
      7651 ,    // 6304
      7651 ,    // 6305
      7652 ,    // 6306
      7652 ,    // 6307
      7653 ,    // 6308
      7654 ,    // 6309
      7654 ,    // 6310
      7655 ,    // 6311
      7655 ,    // 6312
      7656 ,    // 6313
      7656 ,    // 6314
      7657 ,    // 6315
      7657 ,    // 6316
      7658 ,    // 6317
      7659 ,    // 6318
      7659 ,    // 6319
      7660 ,    // 6320
      7660 ,    // 6321
      7661 ,    // 6322
      7661 ,    // 6323
      7662 ,    // 6324
      7662 ,    // 6325
      7663 ,    // 6326
      7663 ,    // 6327
      7664 ,    // 6328
      7665 ,    // 6329
      7665 ,    // 6330
      7666 ,    // 6331
      7666 ,    // 6332
      7667 ,    // 6333
      7667 ,    // 6334
      7668 ,    // 6335
      7668 ,    // 6336
      7669 ,    // 6337
      7670 ,    // 6338
      7670 ,    // 6339
      7671 ,    // 6340
      7671 ,    // 6341
      7672 ,    // 6342
      7672 ,    // 6343
      7673 ,    // 6344
      7673 ,    // 6345
      7674 ,    // 6346
      7674 ,    // 6347
      7675 ,    // 6348
      7676 ,    // 6349
      7676 ,    // 6350
      7677 ,    // 6351
      7677 ,    // 6352
      7678 ,    // 6353
      7678 ,    // 6354
      7679 ,    // 6355
      7679 ,    // 6356
      7680 ,    // 6357
      7680 ,    // 6358
      7681 ,    // 6359
      7681 ,    // 6360
      7682 ,    // 6361
      7683 ,    // 6362
      7683 ,    // 6363
      7684 ,    // 6364
      7684 ,    // 6365
      7685 ,    // 6366
      7685 ,    // 6367
      7686 ,    // 6368
      7686 ,    // 6369
      7687 ,    // 6370
      7687 ,    // 6371
      7688 ,    // 6372
      7688 ,    // 6373
      7689 ,    // 6374
      7690 ,    // 6375
      7690 ,    // 6376
      7691 ,    // 6377
      7691 ,    // 6378
      7692 ,    // 6379
      7692 ,    // 6380
      7693 ,    // 6381
      7693 ,    // 6382
      7694 ,    // 6383
      7694 ,    // 6384
      7695 ,    // 6385
      7695 ,    // 6386
      7696 ,    // 6387
      7696 ,    // 6388
      7697 ,    // 6389
      7698 ,    // 6390
      7698 ,    // 6391
      7699 ,    // 6392
      7699 ,    // 6393
      7700 ,    // 6394
      7700 ,    // 6395
      7701 ,    // 6396
      7701 ,    // 6397
      7702 ,    // 6398
      7702 ,    // 6399
      7703 ,    // 6400
      7703 ,    // 6401
      7704 ,    // 6402
      7704 ,    // 6403
      7705 ,    // 6404
      7705 ,    // 6405
      7706 ,    // 6406
      7707 ,    // 6407
      7707 ,    // 6408
      7708 ,    // 6409
      7708 ,    // 6410
      7709 ,    // 6411
      7709 ,    // 6412
      7710 ,    // 6413
      7710 ,    // 6414
      7711 ,    // 6415
      7711 ,    // 6416
      7712 ,    // 6417
      7712 ,    // 6418
      7713 ,    // 6419
      7713 ,    // 6420
      7714 ,    // 6421
      7714 ,    // 6422
      7715 ,    // 6423
      7715 ,    // 6424
      7716 ,    // 6425
      7716 ,    // 6426
      7717 ,    // 6427
      7718 ,    // 6428
      7718 ,    // 6429
      7719 ,    // 6430
      7719 ,    // 6431
      7720 ,    // 6432
      7720 ,    // 6433
      7721 ,    // 6434
      7721 ,    // 6435
      7722 ,    // 6436
      7722 ,    // 6437
      7723 ,    // 6438
      7723 ,    // 6439
      7724 ,    // 6440
      7724 ,    // 6441
      7725 ,    // 6442
      7725 ,    // 6443
      7726 ,    // 6444
      7726 ,    // 6445
      7727 ,    // 6446
      7727 ,    // 6447
      7728 ,    // 6448
      7728 ,    // 6449
      7729 ,    // 6450
      7729 ,    // 6451
      7730 ,    // 6452
      7730 ,    // 6453
      7731 ,    // 6454
      7731 ,    // 6455
      7732 ,    // 6456
      7732 ,    // 6457
      7733 ,    // 6458
      7734 ,    // 6459
      7734 ,    // 6460
      7735 ,    // 6461
      7735 ,    // 6462
      7736 ,    // 6463
      7736 ,    // 6464
      7737 ,    // 6465
      7737 ,    // 6466
      7738 ,    // 6467
      7738 ,    // 6468
      7739 ,    // 6469
      7739 ,    // 6470
      7740 ,    // 6471
      7740 ,    // 6472
      7741 ,    // 6473
      7741 ,    // 6474
      7742 ,    // 6475
      7742 ,    // 6476
      7743 ,    // 6477
      7743 ,    // 6478
      7744 ,    // 6479
      7744 ,    // 6480
      7745 ,    // 6481
      7745 ,    // 6482
      7746 ,    // 6483
      7746 ,    // 6484
      7747 ,    // 6485
      7747 ,    // 6486
      7748 ,    // 6487
      7748 ,    // 6488
      7749 ,    // 6489
      7749 ,    // 6490
      7750 ,    // 6491
      7750 ,    // 6492
      7751 ,    // 6493
      7751 ,    // 6494
      7752 ,    // 6495
      7752 ,    // 6496
      7753 ,    // 6497
      7753 ,    // 6498
      7754 ,    // 6499
      7754 ,    // 6500
      7755 ,    // 6501
      7755 ,    // 6502
      7756 ,    // 6503
      7756 ,    // 6504
      7757 ,    // 6505
      7757 ,    // 6506
      7758 ,    // 6507
      7758 ,    // 6508
      7759 ,    // 6509
      7759 ,    // 6510
      7760 ,    // 6511
      7760 ,    // 6512
      7761 ,    // 6513
      7761 ,    // 6514
      7762 ,    // 6515
      7762 ,    // 6516
      7763 ,    // 6517
      7763 ,    // 6518
      7764 ,    // 6519
      7764 ,    // 6520
      7765 ,    // 6521
      7765 ,    // 6522
      7766 ,    // 6523
      7766 ,    // 6524
      7767 ,    // 6525
      7767 ,    // 6526
      7768 ,    // 6527
      7768 ,    // 6528
      7769 ,    // 6529
      7769 ,    // 6530
      7770 ,    // 6531
      7770 ,    // 6532
      7771 ,    // 6533
      7771 ,    // 6534
      7772 ,    // 6535
      7772 ,    // 6536
      7773 ,    // 6537
      7773 ,    // 6538
      7774 ,    // 6539
      7774 ,    // 6540
      7775 ,    // 6541
      7775 ,    // 6542
      7775 ,    // 6543
      7776 ,    // 6544
      7776 ,    // 6545
      7777 ,    // 6546
      7777 ,    // 6547
      7778 ,    // 6548
      7778 ,    // 6549
      7779 ,    // 6550
      7779 ,    // 6551
      7780 ,    // 6552
      7780 ,    // 6553
      7781 ,    // 6554
      7781 ,    // 6555
      7782 ,    // 6556
      7782 ,    // 6557
      7783 ,    // 6558
      7783 ,    // 6559
      7784 ,    // 6560
      7784 ,    // 6561
      7785 ,    // 6562
      7785 ,    // 6563
      7786 ,    // 6564
      7786 ,    // 6565
      7787 ,    // 6566
      7787 ,    // 6567
      7788 ,    // 6568
      7788 ,    // 6569
      7789 ,    // 6570
      7789 ,    // 6571
      7790 ,    // 6572
      7790 ,    // 6573
      7790 ,    // 6574
      7791 ,    // 6575
      7791 ,    // 6576
      7792 ,    // 6577
      7792 ,    // 6578
      7793 ,    // 6579
      7793 ,    // 6580
      7794 ,    // 6581
      7794 ,    // 6582
      7795 ,    // 6583
      7795 ,    // 6584
      7796 ,    // 6585
      7796 ,    // 6586
      7797 ,    // 6587
      7797 ,    // 6588
      7798 ,    // 6589
      7798 ,    // 6590
      7799 ,    // 6591
      7799 ,    // 6592
      7800 ,    // 6593
      7800 ,    // 6594
      7800 ,    // 6595
      7801 ,    // 6596
      7801 ,    // 6597
      7802 ,    // 6598
      7802 ,    // 6599
      7803 ,    // 6600
      7803 ,    // 6601
      7804 ,    // 6602
      7804 ,    // 6603
      7805 ,    // 6604
      7805 ,    // 6605
      7806 ,    // 6606
      7806 ,    // 6607
      7807 ,    // 6608
      7807 ,    // 6609
      7808 ,    // 6610
      7808 ,    // 6611
      7808 ,    // 6612
      7809 ,    // 6613
      7809 ,    // 6614
      7810 ,    // 6615
      7810 ,    // 6616
      7811 ,    // 6617
      7811 ,    // 6618
      7812 ,    // 6619
      7812 ,    // 6620
      7813 ,    // 6621
      7813 ,    // 6622
      7814 ,    // 6623
      7814 ,    // 6624
      7815 ,    // 6625
      7815 ,    // 6626
      7815 ,    // 6627
      7816 ,    // 6628
      7816 ,    // 6629
      7817 ,    // 6630
      7817 ,    // 6631
      7818 ,    // 6632
      7818 ,    // 6633
      7819 ,    // 6634
      7819 ,    // 6635
      7820 ,    // 6636
      7820 ,    // 6637
      7821 ,    // 6638
      7821 ,    // 6639
      7821 ,    // 6640
      7822 ,    // 6641
      7822 ,    // 6642
      7823 ,    // 6643
      7823 ,    // 6644
      7824 ,    // 6645
      7824 ,    // 6646
      7825 ,    // 6647
      7825 ,    // 6648
      7826 ,    // 6649
      7826 ,    // 6650
      7827 ,    // 6651
      7827 ,    // 6652
      7827 ,    // 6653
      7828 ,    // 6654
      7828 ,    // 6655
      7829 ,    // 6656
      7829 ,    // 6657
      7830 ,    // 6658
      7830 ,    // 6659
      7831 ,    // 6660
      7831 ,    // 6661
      7832 ,    // 6662
      7832 ,    // 6663
      7832 ,    // 6664
      7833 ,    // 6665
      7833 ,    // 6666
      7834 ,    // 6667
      7834 ,    // 6668
      7835 ,    // 6669
      7835 ,    // 6670
      7836 ,    // 6671
      7836 ,    // 6672
      7836 ,    // 6673
      7837 ,    // 6674
      7837 ,    // 6675
      7838 ,    // 6676
      7838 ,    // 6677
      7839 ,    // 6678
      7839 ,    // 6679
      7840 ,    // 6680
      7840 ,    // 6681
      7841 ,    // 6682
      7841 ,    // 6683
      7841 ,    // 6684
      7842 ,    // 6685
      7842 ,    // 6686
      7843 ,    // 6687
      7843 ,    // 6688
      7844 ,    // 6689
      7844 ,    // 6690
      7845 ,    // 6691
      7845 ,    // 6692
      7845 ,    // 6693
      7846 ,    // 6694
      7846 ,    // 6695
      7847 ,    // 6696
      7847 ,    // 6697
      7848 ,    // 6698
      7848 ,    // 6699
      7849 ,    // 6700
      7849 ,    // 6701
      7849 ,    // 6702
      7850 ,    // 6703
      7850 ,    // 6704
      7851 ,    // 6705
      7851 ,    // 6706
      7852 ,    // 6707
      7852 ,    // 6708
      7853 ,    // 6709
      7853 ,    // 6710
      7853 ,    // 6711
      7854 ,    // 6712
      7854 ,    // 6713
      7855 ,    // 6714
      7855 ,    // 6715
      7856 ,    // 6716
      7856 ,    // 6717
      7856 ,    // 6718
      7857 ,    // 6719
      7857 ,    // 6720
      7858 ,    // 6721
      7858 ,    // 6722
      7859 ,    // 6723
      7859 ,    // 6724
      7860 ,    // 6725
      7860 ,    // 6726
      7860 ,    // 6727
      7861 ,    // 6728
      7861 ,    // 6729
      7862 ,    // 6730
      7862 ,    // 6731
      7863 ,    // 6732
      7863 ,    // 6733
      7863 ,    // 6734
      7864 ,    // 6735
      7864 ,    // 6736
      7865 ,    // 6737
      7865 ,    // 6738
      7866 ,    // 6739
      7866 ,    // 6740
      7866 ,    // 6741
      7867 ,    // 6742
      7867 ,    // 6743
      7868 ,    // 6744
      7868 ,    // 6745
      7869 ,    // 6746
      7869 ,    // 6747
      7869 ,    // 6748
      7870 ,    // 6749
      7870 ,    // 6750
      7871 ,    // 6751
      7871 ,    // 6752
      7872 ,    // 6753
      7872 ,    // 6754
      7872 ,    // 6755
      7873 ,    // 6756
      7873 ,    // 6757
      7874 ,    // 6758
      7874 ,    // 6759
      7875 ,    // 6760
      7875 ,    // 6761
      7875 ,    // 6762
      7876 ,    // 6763
      7876 ,    // 6764
      7877 ,    // 6765
      7877 ,    // 6766
      7878 ,    // 6767
      7878 ,    // 6768
      7878 ,    // 6769
      7879 ,    // 6770
      7879 ,    // 6771
      7880 ,    // 6772
      7880 ,    // 6773
      7881 ,    // 6774
      7881 ,    // 6775
      7881 ,    // 6776
      7882 ,    // 6777
      7882 ,    // 6778
      7883 ,    // 6779
      7883 ,    // 6780
      7883 ,    // 6781
      7884 ,    // 6782
      7884 ,    // 6783
      7885 ,    // 6784
      7885 ,    // 6785
      7886 ,    // 6786
      7886 ,    // 6787
      7886 ,    // 6788
      7887 ,    // 6789
      7887 ,    // 6790
      7888 ,    // 6791
      7888 ,    // 6792
      7888 ,    // 6793
      7889 ,    // 6794
      7889 ,    // 6795
      7890 ,    // 6796
      7890 ,    // 6797
      7891 ,    // 6798
      7891 ,    // 6799
      7891 ,    // 6800
      7892 ,    // 6801
      7892 ,    // 6802
      7893 ,    // 6803
      7893 ,    // 6804
      7893 ,    // 6805
      7894 ,    // 6806
      7894 ,    // 6807
      7895 ,    // 6808
      7895 ,    // 6809
      7895 ,    // 6810
      7896 ,    // 6811
      7896 ,    // 6812
      7897 ,    // 6813
      7897 ,    // 6814
      7898 ,    // 6815
      7898 ,    // 6816
      7898 ,    // 6817
      7899 ,    // 6818
      7899 ,    // 6819
      7900 ,    // 6820
      7900 ,    // 6821
      7900 ,    // 6822
      7901 ,    // 6823
      7901 ,    // 6824
      7902 ,    // 6825
      7902 ,    // 6826
      7902 ,    // 6827
      7903 ,    // 6828
      7903 ,    // 6829
      7904 ,    // 6830
      7904 ,    // 6831
      7904 ,    // 6832
      7905 ,    // 6833
      7905 ,    // 6834
      7906 ,    // 6835
      7906 ,    // 6836
      7906 ,    // 6837
      7907 ,    // 6838
      7907 ,    // 6839
      7908 ,    // 6840
      7908 ,    // 6841
      7908 ,    // 6842
      7909 ,    // 6843
      7909 ,    // 6844
      7910 ,    // 6845
      7910 ,    // 6846
      7910 ,    // 6847
      7911 ,    // 6848
      7911 ,    // 6849
      7912 ,    // 6850
      7912 ,    // 6851
      7912 ,    // 6852
      7913 ,    // 6853
      7913 ,    // 6854
      7914 ,    // 6855
      7914 ,    // 6856
      7914 ,    // 6857
      7915 ,    // 6858
      7915 ,    // 6859
      7916 ,    // 6860
      7916 ,    // 6861
      7916 ,    // 6862
      7917 ,    // 6863
      7917 ,    // 6864
      7918 ,    // 6865
      7918 ,    // 6866
      7918 ,    // 6867
      7919 ,    // 6868
      7919 ,    // 6869
      7920 ,    // 6870
      7920 ,    // 6871
      7920 ,    // 6872
      7921 ,    // 6873
      7921 ,    // 6874
      7922 ,    // 6875
      7922 ,    // 6876
      7922 ,    // 6877
      7923 ,    // 6878
      7923 ,    // 6879
      7924 ,    // 6880
      7924 ,    // 6881
      7924 ,    // 6882
      7925 ,    // 6883
      7925 ,    // 6884
      7925 ,    // 6885
      7926 ,    // 6886
      7926 ,    // 6887
      7927 ,    // 6888
      7927 ,    // 6889
      7927 ,    // 6890
      7928 ,    // 6891
      7928 ,    // 6892
      7929 ,    // 6893
      7929 ,    // 6894
      7929 ,    // 6895
      7930 ,    // 6896
      7930 ,    // 6897
      7931 ,    // 6898
      7931 ,    // 6899
      7931 ,    // 6900
      7932 ,    // 6901
      7932 ,    // 6902
      7932 ,    // 6903
      7933 ,    // 6904
      7933 ,    // 6905
      7934 ,    // 6906
      7934 ,    // 6907
      7934 ,    // 6908
      7935 ,    // 6909
      7935 ,    // 6910
      7936 ,    // 6911
      7936 ,    // 6912
      7936 ,    // 6913
      7937 ,    // 6914
      7937 ,    // 6915
      7937 ,    // 6916
      7938 ,    // 6917
      7938 ,    // 6918
      7939 ,    // 6919
      7939 ,    // 6920
      7939 ,    // 6921
      7940 ,    // 6922
      7940 ,    // 6923
      7940 ,    // 6924
      7941 ,    // 6925
      7941 ,    // 6926
      7942 ,    // 6927
      7942 ,    // 6928
      7942 ,    // 6929
      7943 ,    // 6930
      7943 ,    // 6931
      7943 ,    // 6932
      7944 ,    // 6933
      7944 ,    // 6934
      7945 ,    // 6935
      7945 ,    // 6936
      7945 ,    // 6937
      7946 ,    // 6938
      7946 ,    // 6939
      7946 ,    // 6940
      7947 ,    // 6941
      7947 ,    // 6942
      7948 ,    // 6943
      7948 ,    // 6944
      7948 ,    // 6945
      7949 ,    // 6946
      7949 ,    // 6947
      7949 ,    // 6948
      7950 ,    // 6949
      7950 ,    // 6950
      7951 ,    // 6951
      7951 ,    // 6952
      7951 ,    // 6953
      7952 ,    // 6954
      7952 ,    // 6955
      7952 ,    // 6956
      7953 ,    // 6957
      7953 ,    // 6958
      7953 ,    // 6959
      7954 ,    // 6960
      7954 ,    // 6961
      7955 ,    // 6962
      7955 ,    // 6963
      7955 ,    // 6964
      7956 ,    // 6965
      7956 ,    // 6966
      7956 ,    // 6967
      7957 ,    // 6968
      7957 ,    // 6969
      7958 ,    // 6970
      7958 ,    // 6971
      7958 ,    // 6972
      7959 ,    // 6973
      7959 ,    // 6974
      7959 ,    // 6975
      7960 ,    // 6976
      7960 ,    // 6977
      7960 ,    // 6978
      7961 ,    // 6979
      7961 ,    // 6980
      7961 ,    // 6981
      7962 ,    // 6982
      7962 ,    // 6983
      7963 ,    // 6984
      7963 ,    // 6985
      7963 ,    // 6986
      7964 ,    // 6987
      7964 ,    // 6988
      7964 ,    // 6989
      7965 ,    // 6990
      7965 ,    // 6991
      7965 ,    // 6992
      7966 ,    // 6993
      7966 ,    // 6994
      7967 ,    // 6995
      7967 ,    // 6996
      7967 ,    // 6997
      7968 ,    // 6998
      7968 ,    // 6999
      7968 ,    // 7000
      7969 ,    // 7001
      7969 ,    // 7002
      7969 ,    // 7003
      7970 ,    // 7004
      7970 ,    // 7005
      7970 ,    // 7006
      7971 ,    // 7007
      7971 ,    // 7008
      7971 ,    // 7009
      7972 ,    // 7010
      7972 ,    // 7011
      7973 ,    // 7012
      7973 ,    // 7013
      7973 ,    // 7014
      7974 ,    // 7015
      7974 ,    // 7016
      7974 ,    // 7017
      7975 ,    // 7018
      7975 ,    // 7019
      7975 ,    // 7020
      7976 ,    // 7021
      7976 ,    // 7022
      7976 ,    // 7023
      7977 ,    // 7024
      7977 ,    // 7025
      7977 ,    // 7026
      7978 ,    // 7027
      7978 ,    // 7028
      7978 ,    // 7029
      7979 ,    // 7030
      7979 ,    // 7031
      7980 ,    // 7032
      7980 ,    // 7033
      7980 ,    // 7034
      7981 ,    // 7035
      7981 ,    // 7036
      7981 ,    // 7037
      7982 ,    // 7038
      7982 ,    // 7039
      7982 ,    // 7040
      7983 ,    // 7041
      7983 ,    // 7042
      7983 ,    // 7043
      7984 ,    // 7044
      7984 ,    // 7045
      7984 ,    // 7046
      7985 ,    // 7047
      7985 ,    // 7048
      7985 ,    // 7049
      7986 ,    // 7050
      7986 ,    // 7051
      7986 ,    // 7052
      7987 ,    // 7053
      7987 ,    // 7054
      7987 ,    // 7055
      7988 ,    // 7056
      7988 ,    // 7057
      7988 ,    // 7058
      7989 ,    // 7059
      7989 ,    // 7060
      7989 ,    // 7061
      7990 ,    // 7062
      7990 ,    // 7063
      7990 ,    // 7064
      7991 ,    // 7065
      7991 ,    // 7066
      7991 ,    // 7067
      7992 ,    // 7068
      7992 ,    // 7069
      7992 ,    // 7070
      7993 ,    // 7071
      7993 ,    // 7072
      7993 ,    // 7073
      7994 ,    // 7074
      7994 ,    // 7075
      7994 ,    // 7076
      7995 ,    // 7077
      7995 ,    // 7078
      7995 ,    // 7079
      7996 ,    // 7080
      7996 ,    // 7081
      7996 ,    // 7082
      7997 ,    // 7083
      7997 ,    // 7084
      7997 ,    // 7085
      7998 ,    // 7086
      7998 ,    // 7087
      7998 ,    // 7088
      7999 ,    // 7089
      7999 ,    // 7090
      7999 ,    // 7091
      8000 ,    // 7092
      8000 ,    // 7093
      8000 ,    // 7094
      8001 ,    // 7095
      8001 ,    // 7096
      8001 ,    // 7097
      8002 ,    // 7098
      8002 ,    // 7099
      8002 ,    // 7100
      8003 ,    // 7101
      8003 ,    // 7102
      8003 ,    // 7103
      8004 ,    // 7104
      8004 ,    // 7105
      8004 ,    // 7106
      8005 ,    // 7107
      8005 ,    // 7108
      8005 ,    // 7109
      8006 ,    // 7110
      8006 ,    // 7111
      8006 ,    // 7112
      8007 ,    // 7113
      8007 ,    // 7114
      8007 ,    // 7115
      8008 ,    // 7116
      8008 ,    // 7117
      8008 ,    // 7118
      8009 ,    // 7119
      8009 ,    // 7120
      8009 ,    // 7121
      8009 ,    // 7122
      8010 ,    // 7123
      8010 ,    // 7124
      8010 ,    // 7125
      8011 ,    // 7126
      8011 ,    // 7127
      8011 ,    // 7128
      8012 ,    // 7129
      8012 ,    // 7130
      8012 ,    // 7131
      8013 ,    // 7132
      8013 ,    // 7133
      8013 ,    // 7134
      8014 ,    // 7135
      8014 ,    // 7136
      8014 ,    // 7137
      8015 ,    // 7138
      8015 ,    // 7139
      8015 ,    // 7140
      8015 ,    // 7141
      8016 ,    // 7142
      8016 ,    // 7143
      8016 ,    // 7144
      8017 ,    // 7145
      8017 ,    // 7146
      8017 ,    // 7147
      8018 ,    // 7148
      8018 ,    // 7149
      8018 ,    // 7150
      8019 ,    // 7151
      8019 ,    // 7152
      8019 ,    // 7153
      8020 ,    // 7154
      8020 ,    // 7155
      8020 ,    // 7156
      8020 ,    // 7157
      8021 ,    // 7158
      8021 ,    // 7159
      8021 ,    // 7160
      8022 ,    // 7161
      8022 ,    // 7162
      8022 ,    // 7163
      8023 ,    // 7164
      8023 ,    // 7165
      8023 ,    // 7166
      8024 ,    // 7167
      8024 ,    // 7168
      8024 ,    // 7169
      8024 ,    // 7170
      8025 ,    // 7171
      8025 ,    // 7172
      8025 ,    // 7173
      8026 ,    // 7174
      8026 ,    // 7175
      8026 ,    // 7176
      8027 ,    // 7177
      8027 ,    // 7178
      8027 ,    // 7179
      8028 ,    // 7180
      8028 ,    // 7181
      8028 ,    // 7182
      8028 ,    // 7183
      8029 ,    // 7184
      8029 ,    // 7185
      8029 ,    // 7186
      8030 ,    // 7187
      8030 ,    // 7188
      8030 ,    // 7189
      8031 ,    // 7190
      8031 ,    // 7191
      8031 ,    // 7192
      8031 ,    // 7193
      8032 ,    // 7194
      8032 ,    // 7195
      8032 ,    // 7196
      8033 ,    // 7197
      8033 ,    // 7198
      8033 ,    // 7199
      8034 ,    // 7200
      8034 ,    // 7201
      8034 ,    // 7202
      8034 ,    // 7203
      8035 ,    // 7204
      8035 ,    // 7205
      8035 ,    // 7206
      8036 ,    // 7207
      8036 ,    // 7208
      8036 ,    // 7209
      8036 ,    // 7210
      8037 ,    // 7211
      8037 ,    // 7212
      8037 ,    // 7213
      8038 ,    // 7214
      8038 ,    // 7215
      8038 ,    // 7216
      8039 ,    // 7217
      8039 ,    // 7218
      8039 ,    // 7219
      8039 ,    // 7220
      8040 ,    // 7221
      8040 ,    // 7222
      8040 ,    // 7223
      8041 ,    // 7224
      8041 ,    // 7225
      8041 ,    // 7226
      8041 ,    // 7227
      8042 ,    // 7228
      8042 ,    // 7229
      8042 ,    // 7230
      8043 ,    // 7231
      8043 ,    // 7232
      8043 ,    // 7233
      8043 ,    // 7234
      8044 ,    // 7235
      8044 ,    // 7236
      8044 ,    // 7237
      8045 ,    // 7238
      8045 ,    // 7239
      8045 ,    // 7240
      8045 ,    // 7241
      8046 ,    // 7242
      8046 ,    // 7243
      8046 ,    // 7244
      8047 ,    // 7245
      8047 ,    // 7246
      8047 ,    // 7247
      8047 ,    // 7248
      8048 ,    // 7249
      8048 ,    // 7250
      8048 ,    // 7251
      8049 ,    // 7252
      8049 ,    // 7253
      8049 ,    // 7254
      8049 ,    // 7255
      8050 ,    // 7256
      8050 ,    // 7257
      8050 ,    // 7258
      8050 ,    // 7259
      8051 ,    // 7260
      8051 ,    // 7261
      8051 ,    // 7262
      8052 ,    // 7263
      8052 ,    // 7264
      8052 ,    // 7265
      8052 ,    // 7266
      8053 ,    // 7267
      8053 ,    // 7268
      8053 ,    // 7269
      8054 ,    // 7270
      8054 ,    // 7271
      8054 ,    // 7272
      8054 ,    // 7273
      8055 ,    // 7274
      8055 ,    // 7275
      8055 ,    // 7276
      8055 ,    // 7277
      8056 ,    // 7278
      8056 ,    // 7279
      8056 ,    // 7280
      8057 ,    // 7281
      8057 ,    // 7282
      8057 ,    // 7283
      8057 ,    // 7284
      8058 ,    // 7285
      8058 ,    // 7286
      8058 ,    // 7287
      8058 ,    // 7288
      8059 ,    // 7289
      8059 ,    // 7290
      8059 ,    // 7291
      8060 ,    // 7292
      8060 ,    // 7293
      8060 ,    // 7294
      8060 ,    // 7295
      8061 ,    // 7296
      8061 ,    // 7297
      8061 ,    // 7298
      8061 ,    // 7299
      8062 ,    // 7300
      8062 ,    // 7301
      8062 ,    // 7302
      8062 ,    // 7303
      8063 ,    // 7304
      8063 ,    // 7305
      8063 ,    // 7306
      8064 ,    // 7307
      8064 ,    // 7308
      8064 ,    // 7309
      8064 ,    // 7310
      8065 ,    // 7311
      8065 ,    // 7312
      8065 ,    // 7313
      8065 ,    // 7314
      8066 ,    // 7315
      8066 ,    // 7316
      8066 ,    // 7317
      8066 ,    // 7318
      8067 ,    // 7319
      8067 ,    // 7320
      8067 ,    // 7321
      8067 ,    // 7322
      8068 ,    // 7323
      8068 ,    // 7324
      8068 ,    // 7325
      8069 ,    // 7326
      8069 ,    // 7327
      8069 ,    // 7328
      8069 ,    // 7329
      8070 ,    // 7330
      8070 ,    // 7331
      8070 ,    // 7332
      8070 ,    // 7333
      8071 ,    // 7334
      8071 ,    // 7335
      8071 ,    // 7336
      8071 ,    // 7337
      8072 ,    // 7338
      8072 ,    // 7339
      8072 ,    // 7340
      8072 ,    // 7341
      8073 ,    // 7342
      8073 ,    // 7343
      8073 ,    // 7344
      8073 ,    // 7345
      8074 ,    // 7346
      8074 ,    // 7347
      8074 ,    // 7348
      8074 ,    // 7349
      8075 ,    // 7350
      8075 ,    // 7351
      8075 ,    // 7352
      8075 ,    // 7353
      8076 ,    // 7354
      8076 ,    // 7355
      8076 ,    // 7356
      8076 ,    // 7357
      8077 ,    // 7358
      8077 ,    // 7359
      8077 ,    // 7360
      8077 ,    // 7361
      8078 ,    // 7362
      8078 ,    // 7363
      8078 ,    // 7364
      8078 ,    // 7365
      8079 ,    // 7366
      8079 ,    // 7367
      8079 ,    // 7368
      8079 ,    // 7369
      8080 ,    // 7370
      8080 ,    // 7371
      8080 ,    // 7372
      8080 ,    // 7373
      8081 ,    // 7374
      8081 ,    // 7375
      8081 ,    // 7376
      8081 ,    // 7377
      8082 ,    // 7378
      8082 ,    // 7379
      8082 ,    // 7380
      8082 ,    // 7381
      8083 ,    // 7382
      8083 ,    // 7383
      8083 ,    // 7384
      8083 ,    // 7385
      8084 ,    // 7386
      8084 ,    // 7387
      8084 ,    // 7388
      8084 ,    // 7389
      8085 ,    // 7390
      8085 ,    // 7391
      8085 ,    // 7392
      8085 ,    // 7393
      8085 ,    // 7394
      8086 ,    // 7395
      8086 ,    // 7396
      8086 ,    // 7397
      8086 ,    // 7398
      8087 ,    // 7399
      8087 ,    // 7400
      8087 ,    // 7401
      8087 ,    // 7402
      8088 ,    // 7403
      8088 ,    // 7404
      8088 ,    // 7405
      8088 ,    // 7406
      8089 ,    // 7407
      8089 ,    // 7408
      8089 ,    // 7409
      8089 ,    // 7410
      8089 ,    // 7411
      8090 ,    // 7412
      8090 ,    // 7413
      8090 ,    // 7414
      8090 ,    // 7415
      8091 ,    // 7416
      8091 ,    // 7417
      8091 ,    // 7418
      8091 ,    // 7419
      8092 ,    // 7420
      8092 ,    // 7421
      8092 ,    // 7422
      8092 ,    // 7423
      8093 ,    // 7424
      8093 ,    // 7425
      8093 ,    // 7426
      8093 ,    // 7427
      8093 ,    // 7428
      8094 ,    // 7429
      8094 ,    // 7430
      8094 ,    // 7431
      8094 ,    // 7432
      8095 ,    // 7433
      8095 ,    // 7434
      8095 ,    // 7435
      8095 ,    // 7436
      8095 ,    // 7437
      8096 ,    // 7438
      8096 ,    // 7439
      8096 ,    // 7440
      8096 ,    // 7441
      8097 ,    // 7442
      8097 ,    // 7443
      8097 ,    // 7444
      8097 ,    // 7445
      8098 ,    // 7446
      8098 ,    // 7447
      8098 ,    // 7448
      8098 ,    // 7449
      8098 ,    // 7450
      8099 ,    // 7451
      8099 ,    // 7452
      8099 ,    // 7453
      8099 ,    // 7454
      8100 ,    // 7455
      8100 ,    // 7456
      8100 ,    // 7457
      8100 ,    // 7458
      8100 ,    // 7459
      8101 ,    // 7460
      8101 ,    // 7461
      8101 ,    // 7462
      8101 ,    // 7463
      8101 ,    // 7464
      8102 ,    // 7465
      8102 ,    // 7466
      8102 ,    // 7467
      8102 ,    // 7468
      8103 ,    // 7469
      8103 ,    // 7470
      8103 ,    // 7471
      8103 ,    // 7472
      8103 ,    // 7473
      8104 ,    // 7474
      8104 ,    // 7475
      8104 ,    // 7476
      8104 ,    // 7477
      8105 ,    // 7478
      8105 ,    // 7479
      8105 ,    // 7480
      8105 ,    // 7481
      8105 ,    // 7482
      8106 ,    // 7483
      8106 ,    // 7484
      8106 ,    // 7485
      8106 ,    // 7486
      8106 ,    // 7487
      8107 ,    // 7488
      8107 ,    // 7489
      8107 ,    // 7490
      8107 ,    // 7491
      8107 ,    // 7492
      8108 ,    // 7493
      8108 ,    // 7494
      8108 ,    // 7495
      8108 ,    // 7496
      8109 ,    // 7497
      8109 ,    // 7498
      8109 ,    // 7499
      8109 ,    // 7500
      8109 ,    // 7501
      8110 ,    // 7502
      8110 ,    // 7503
      8110 ,    // 7504
      8110 ,    // 7505
      8110 ,    // 7506
      8111 ,    // 7507
      8111 ,    // 7508
      8111 ,    // 7509
      8111 ,    // 7510
      8111 ,    // 7511
      8112 ,    // 7512
      8112 ,    // 7513
      8112 ,    // 7514
      8112 ,    // 7515
      8112 ,    // 7516
      8113 ,    // 7517
      8113 ,    // 7518
      8113 ,    // 7519
      8113 ,    // 7520
      8113 ,    // 7521
      8114 ,    // 7522
      8114 ,    // 7523
      8114 ,    // 7524
      8114 ,    // 7525
      8114 ,    // 7526
      8115 ,    // 7527
      8115 ,    // 7528
      8115 ,    // 7529
      8115 ,    // 7530
      8115 ,    // 7531
      8116 ,    // 7532
      8116 ,    // 7533
      8116 ,    // 7534
      8116 ,    // 7535
      8116 ,    // 7536
      8117 ,    // 7537
      8117 ,    // 7538
      8117 ,    // 7539
      8117 ,    // 7540
      8117 ,    // 7541
      8118 ,    // 7542
      8118 ,    // 7543
      8118 ,    // 7544
      8118 ,    // 7545
      8118 ,    // 7546
      8119 ,    // 7547
      8119 ,    // 7548
      8119 ,    // 7549
      8119 ,    // 7550
      8119 ,    // 7551
      8120 ,    // 7552
      8120 ,    // 7553
      8120 ,    // 7554
      8120 ,    // 7555
      8120 ,    // 7556
      8120 ,    // 7557
      8121 ,    // 7558
      8121 ,    // 7559
      8121 ,    // 7560
      8121 ,    // 7561
      8121 ,    // 7562
      8122 ,    // 7563
      8122 ,    // 7564
      8122 ,    // 7565
      8122 ,    // 7566
      8122 ,    // 7567
      8123 ,    // 7568
      8123 ,    // 7569
      8123 ,    // 7570
      8123 ,    // 7571
      8123 ,    // 7572
      8124 ,    // 7573
      8124 ,    // 7574
      8124 ,    // 7575
      8124 ,    // 7576
      8124 ,    // 7577
      8124 ,    // 7578
      8125 ,    // 7579
      8125 ,    // 7580
      8125 ,    // 7581
      8125 ,    // 7582
      8125 ,    // 7583
      8126 ,    // 7584
      8126 ,    // 7585
      8126 ,    // 7586
      8126 ,    // 7587
      8126 ,    // 7588
      8126 ,    // 7589
      8127 ,    // 7590
      8127 ,    // 7591
      8127 ,    // 7592
      8127 ,    // 7593
      8127 ,    // 7594
      8128 ,    // 7595
      8128 ,    // 7596
      8128 ,    // 7597
      8128 ,    // 7598
      8128 ,    // 7599
      8128 ,    // 7600
      8129 ,    // 7601
      8129 ,    // 7602
      8129 ,    // 7603
      8129 ,    // 7604
      8129 ,    // 7605
      8129 ,    // 7606
      8130 ,    // 7607
      8130 ,    // 7608
      8130 ,    // 7609
      8130 ,    // 7610
      8130 ,    // 7611
      8131 ,    // 7612
      8131 ,    // 7613
      8131 ,    // 7614
      8131 ,    // 7615
      8131 ,    // 7616
      8131 ,    // 7617
      8132 ,    // 7618
      8132 ,    // 7619
      8132 ,    // 7620
      8132 ,    // 7621
      8132 ,    // 7622
      8132 ,    // 7623
      8133 ,    // 7624
      8133 ,    // 7625
      8133 ,    // 7626
      8133 ,    // 7627
      8133 ,    // 7628
      8133 ,    // 7629
      8134 ,    // 7630
      8134 ,    // 7631
      8134 ,    // 7632
      8134 ,    // 7633
      8134 ,    // 7634
      8134 ,    // 7635
      8135 ,    // 7636
      8135 ,    // 7637
      8135 ,    // 7638
      8135 ,    // 7639
      8135 ,    // 7640
      8135 ,    // 7641
      8136 ,    // 7642
      8136 ,    // 7643
      8136 ,    // 7644
      8136 ,    // 7645
      8136 ,    // 7646
      8136 ,    // 7647
      8137 ,    // 7648
      8137 ,    // 7649
      8137 ,    // 7650
      8137 ,    // 7651
      8137 ,    // 7652
      8137 ,    // 7653
      8138 ,    // 7654
      8138 ,    // 7655
      8138 ,    // 7656
      8138 ,    // 7657
      8138 ,    // 7658
      8138 ,    // 7659
      8139 ,    // 7660
      8139 ,    // 7661
      8139 ,    // 7662
      8139 ,    // 7663
      8139 ,    // 7664
      8139 ,    // 7665
      8139 ,    // 7666
      8140 ,    // 7667
      8140 ,    // 7668
      8140 ,    // 7669
      8140 ,    // 7670
      8140 ,    // 7671
      8140 ,    // 7672
      8141 ,    // 7673
      8141 ,    // 7674
      8141 ,    // 7675
      8141 ,    // 7676
      8141 ,    // 7677
      8141 ,    // 7678
      8142 ,    // 7679
      8142 ,    // 7680
      8142 ,    // 7681
      8142 ,    // 7682
      8142 ,    // 7683
      8142 ,    // 7684
      8142 ,    // 7685
      8143 ,    // 7686
      8143 ,    // 7687
      8143 ,    // 7688
      8143 ,    // 7689
      8143 ,    // 7690
      8143 ,    // 7691
      8143 ,    // 7692
      8144 ,    // 7693
      8144 ,    // 7694
      8144 ,    // 7695
      8144 ,    // 7696
      8144 ,    // 7697
      8144 ,    // 7698
      8145 ,    // 7699
      8145 ,    // 7700
      8145 ,    // 7701
      8145 ,    // 7702
      8145 ,    // 7703
      8145 ,    // 7704
      8145 ,    // 7705
      8146 ,    // 7706
      8146 ,    // 7707
      8146 ,    // 7708
      8146 ,    // 7709
      8146 ,    // 7710
      8146 ,    // 7711
      8146 ,    // 7712
      8147 ,    // 7713
      8147 ,    // 7714
      8147 ,    // 7715
      8147 ,    // 7716
      8147 ,    // 7717
      8147 ,    // 7718
      8147 ,    // 7719
      8148 ,    // 7720
      8148 ,    // 7721
      8148 ,    // 7722
      8148 ,    // 7723
      8148 ,    // 7724
      8148 ,    // 7725
      8148 ,    // 7726
      8149 ,    // 7727
      8149 ,    // 7728
      8149 ,    // 7729
      8149 ,    // 7730
      8149 ,    // 7731
      8149 ,    // 7732
      8149 ,    // 7733
      8150 ,    // 7734
      8150 ,    // 7735
      8150 ,    // 7736
      8150 ,    // 7737
      8150 ,    // 7738
      8150 ,    // 7739
      8150 ,    // 7740
      8150 ,    // 7741
      8151 ,    // 7742
      8151 ,    // 7743
      8151 ,    // 7744
      8151 ,    // 7745
      8151 ,    // 7746
      8151 ,    // 7747
      8151 ,    // 7748
      8152 ,    // 7749
      8152 ,    // 7750
      8152 ,    // 7751
      8152 ,    // 7752
      8152 ,    // 7753
      8152 ,    // 7754
      8152 ,    // 7755
      8152 ,    // 7756
      8153 ,    // 7757
      8153 ,    // 7758
      8153 ,    // 7759
      8153 ,    // 7760
      8153 ,    // 7761
      8153 ,    // 7762
      8153 ,    // 7763
      8154 ,    // 7764
      8154 ,    // 7765
      8154 ,    // 7766
      8154 ,    // 7767
      8154 ,    // 7768
      8154 ,    // 7769
      8154 ,    // 7770
      8154 ,    // 7771
      8155 ,    // 7772
      8155 ,    // 7773
      8155 ,    // 7774
      8155 ,    // 7775
      8155 ,    // 7776
      8155 ,    // 7777
      8155 ,    // 7778
      8155 ,    // 7779
      8156 ,    // 7780
      8156 ,    // 7781
      8156 ,    // 7782
      8156 ,    // 7783
      8156 ,    // 7784
      8156 ,    // 7785
      8156 ,    // 7786
      8156 ,    // 7787
      8157 ,    // 7788
      8157 ,    // 7789
      8157 ,    // 7790
      8157 ,    // 7791
      8157 ,    // 7792
      8157 ,    // 7793
      8157 ,    // 7794
      8157 ,    // 7795
      8157 ,    // 7796
      8158 ,    // 7797
      8158 ,    // 7798
      8158 ,    // 7799
      8158 ,    // 7800
      8158 ,    // 7801
      8158 ,    // 7802
      8158 ,    // 7803
      8158 ,    // 7804
      8159 ,    // 7805
      8159 ,    // 7806
      8159 ,    // 7807
      8159 ,    // 7808
      8159 ,    // 7809
      8159 ,    // 7810
      8159 ,    // 7811
      8159 ,    // 7812
      8159 ,    // 7813
      8160 ,    // 7814
      8160 ,    // 7815
      8160 ,    // 7816
      8160 ,    // 7817
      8160 ,    // 7818
      8160 ,    // 7819
      8160 ,    // 7820
      8160 ,    // 7821
      8160 ,    // 7822
      8161 ,    // 7823
      8161 ,    // 7824
      8161 ,    // 7825
      8161 ,    // 7826
      8161 ,    // 7827
      8161 ,    // 7828
      8161 ,    // 7829
      8161 ,    // 7830
      8161 ,    // 7831
      8162 ,    // 7832
      8162 ,    // 7833
      8162 ,    // 7834
      8162 ,    // 7835
      8162 ,    // 7836
      8162 ,    // 7837
      8162 ,    // 7838
      8162 ,    // 7839
      8162 ,    // 7840
      8163 ,    // 7841
      8163 ,    // 7842
      8163 ,    // 7843
      8163 ,    // 7844
      8163 ,    // 7845
      8163 ,    // 7846
      8163 ,    // 7847
      8163 ,    // 7848
      8163 ,    // 7849
      8163 ,    // 7850
      8164 ,    // 7851
      8164 ,    // 7852
      8164 ,    // 7853
      8164 ,    // 7854
      8164 ,    // 7855
      8164 ,    // 7856
      8164 ,    // 7857
      8164 ,    // 7858
      8164 ,    // 7859
      8164 ,    // 7860
      8165 ,    // 7861
      8165 ,    // 7862
      8165 ,    // 7863
      8165 ,    // 7864
      8165 ,    // 7865
      8165 ,    // 7866
      8165 ,    // 7867
      8165 ,    // 7868
      8165 ,    // 7869
      8165 ,    // 7870
      8166 ,    // 7871
      8166 ,    // 7872
      8166 ,    // 7873
      8166 ,    // 7874
      8166 ,    // 7875
      8166 ,    // 7876
      8166 ,    // 7877
      8166 ,    // 7878
      8166 ,    // 7879
      8166 ,    // 7880
      8167 ,    // 7881
      8167 ,    // 7882
      8167 ,    // 7883
      8167 ,    // 7884
      8167 ,    // 7885
      8167 ,    // 7886
      8167 ,    // 7887
      8167 ,    // 7888
      8167 ,    // 7889
      8167 ,    // 7890
      8167 ,    // 7891
      8168 ,    // 7892
      8168 ,    // 7893
      8168 ,    // 7894
      8168 ,    // 7895
      8168 ,    // 7896
      8168 ,    // 7897
      8168 ,    // 7898
      8168 ,    // 7899
      8168 ,    // 7900
      8168 ,    // 7901
      8168 ,    // 7902
      8169 ,    // 7903
      8169 ,    // 7904
      8169 ,    // 7905
      8169 ,    // 7906
      8169 ,    // 7907
      8169 ,    // 7908
      8169 ,    // 7909
      8169 ,    // 7910
      8169 ,    // 7911
      8169 ,    // 7912
      8169 ,    // 7913
      8169 ,    // 7914
      8170 ,    // 7915
      8170 ,    // 7916
      8170 ,    // 7917
      8170 ,    // 7918
      8170 ,    // 7919
      8170 ,    // 7920
      8170 ,    // 7921
      8170 ,    // 7922
      8170 ,    // 7923
      8170 ,    // 7924
      8170 ,    // 7925
      8170 ,    // 7926
      8171 ,    // 7927
      8171 ,    // 7928
      8171 ,    // 7929
      8171 ,    // 7930
      8171 ,    // 7931
      8171 ,    // 7932
      8171 ,    // 7933
      8171 ,    // 7934
      8171 ,    // 7935
      8171 ,    // 7936
      8171 ,    // 7937
      8171 ,    // 7938
      8171 ,    // 7939
      8172 ,    // 7940
      8172 ,    // 7941
      8172 ,    // 7942
      8172 ,    // 7943
      8172 ,    // 7944
      8172 ,    // 7945
      8172 ,    // 7946
      8172 ,    // 7947
      8172 ,    // 7948
      8172 ,    // 7949
      8172 ,    // 7950
      8172 ,    // 7951
      8172 ,    // 7952
      8172 ,    // 7953
      8173 ,    // 7954
      8173 ,    // 7955
      8173 ,    // 7956
      8173 ,    // 7957
      8173 ,    // 7958
      8173 ,    // 7959
      8173 ,    // 7960
      8173 ,    // 7961
      8173 ,    // 7962
      8173 ,    // 7963
      8173 ,    // 7964
      8173 ,    // 7965
      8173 ,    // 7966
      8173 ,    // 7967
      8174 ,    // 7968
      8174 ,    // 7969
      8174 ,    // 7970
      8174 ,    // 7971
      8174 ,    // 7972
      8174 ,    // 7973
      8174 ,    // 7974
      8174 ,    // 7975
      8174 ,    // 7976
      8174 ,    // 7977
      8174 ,    // 7978
      8174 ,    // 7979
      8174 ,    // 7980
      8174 ,    // 7981
      8174 ,    // 7982
      8174 ,    // 7983
      8175 ,    // 7984
      8175 ,    // 7985
      8175 ,    // 7986
      8175 ,    // 7987
      8175 ,    // 7988
      8175 ,    // 7989
      8175 ,    // 7990
      8175 ,    // 7991
      8175 ,    // 7992
      8175 ,    // 7993
      8175 ,    // 7994
      8175 ,    // 7995
      8175 ,    // 7996
      8175 ,    // 7997
      8175 ,    // 7998
      8175 ,    // 7999
      8176 ,    // 8000
      8176 ,    // 8001
      8176 ,    // 8002
      8176 ,    // 8003
      8176 ,    // 8004
      8176 ,    // 8005
      8176 ,    // 8006
      8176 ,    // 8007
      8176 ,    // 8008
      8176 ,    // 8009
      8176 ,    // 8010
      8176 ,    // 8011
      8176 ,    // 8012
      8176 ,    // 8013
      8176 ,    // 8014
      8176 ,    // 8015
      8176 ,    // 8016
      8176 ,    // 8017
      8177 ,    // 8018
      8177 ,    // 8019
      8177 ,    // 8020
      8177 ,    // 8021
      8177 ,    // 8022
      8177 ,    // 8023
      8177 ,    // 8024
      8177 ,    // 8025
      8177 ,    // 8026
      8177 ,    // 8027
      8177 ,    // 8028
      8177 ,    // 8029
      8177 ,    // 8030
      8177 ,    // 8031
      8177 ,    // 8032
      8177 ,    // 8033
      8177 ,    // 8034
      8177 ,    // 8035
      8177 ,    // 8036
      8177 ,    // 8037
      8177 ,    // 8038
      8178 ,    // 8039
      8178 ,    // 8040
      8178 ,    // 8041
      8178 ,    // 8042
      8178 ,    // 8043
      8178 ,    // 8044
      8178 ,    // 8045
      8178 ,    // 8046
      8178 ,    // 8047
      8178 ,    // 8048
      8178 ,    // 8049
      8178 ,    // 8050
      8178 ,    // 8051
      8178 ,    // 8052
      8178 ,    // 8053
      8178 ,    // 8054
      8178 ,    // 8055
      8178 ,    // 8056
      8178 ,    // 8057
      8178 ,    // 8058
      8178 ,    // 8059
      8178 ,    // 8060
      8178 ,    // 8061
      8179 ,    // 8062
      8179 ,    // 8063
      8179 ,    // 8064
      8179 ,    // 8065
      8179 ,    // 8066
      8179 ,    // 8067
      8179 ,    // 8068
      8179 ,    // 8069
      8179 ,    // 8070
      8179 ,    // 8071
      8179 ,    // 8072
      8179 ,    // 8073
      8179 ,    // 8074
      8179 ,    // 8075
      8179 ,    // 8076
      8179 ,    // 8077
      8179 ,    // 8078
      8179 ,    // 8079
      8179 ,    // 8080
      8179 ,    // 8081
      8179 ,    // 8082
      8179 ,    // 8083
      8179 ,    // 8084
      8179 ,    // 8085
      8179 ,    // 8086
      8179 ,    // 8087
      8179 ,    // 8088
      8179 ,    // 8089
      8179 ,    // 8090
      8180 ,    // 8091
      8180 ,    // 8092
      8180 ,    // 8093
      8180 ,    // 8094
      8180 ,    // 8095
      8180 ,    // 8096
      8180 ,    // 8097
      8180 ,    // 8098
      8180 ,    // 8099
      8180 ,    // 8100
      8180 ,    // 8101
      8180 ,    // 8102
      8180 ,    // 8103
      8180 ,    // 8104
      8180 ,    // 8105
      8180 ,    // 8106
      8180 ,    // 8107
      8180 ,    // 8108
      8180 ,    // 8109
      8180 ,    // 8110
      8180 ,    // 8111
      8180 ,    // 8112
      8180 ,    // 8113
      8180 ,    // 8114
      8180 ,    // 8115
      8180 ,    // 8116
      8180 ,    // 8117
      8180 ,    // 8118
      8180 ,    // 8119
      8180 ,    // 8120
      8180 ,    // 8121
      8180 ,    // 8122
      8180 ,    // 8123
      8180 ,    // 8124
      8180 ,    // 8125
      8180 ,    // 8126
      8180 ,    // 8127
      8180 ,    // 8128
      8180 ,    // 8129
      8180 ,    // 8130
      8181 ,    // 8131
      8181 ,    // 8132
      8181 ,    // 8133
      8181 ,    // 8134
      8181 ,    // 8135
      8181 ,    // 8136
      8181 ,    // 8137
      8181 ,    // 8138
      8181 ,    // 8139
      8181 ,    // 8140
      8181 ,    // 8141
      8181 ,    // 8142
      8181 ,    // 8143
      8181 ,    // 8144
      8181 ,    // 8145
      8181 ,    // 8146
      8181 ,    // 8147
      8181 ,    // 8148
      8181 ,    // 8149
      8181 ,    // 8150
      8181 ,    // 8151
      8181 ,    // 8152
      8181 ,    // 8153
      8181 ,    // 8154
      8181 ,    // 8155
      8181 ,    // 8156
      8181 ,    // 8157
      8181 ,    // 8158
      8181 ,    // 8159
      8181 ,    // 8160
      8181 ,    // 8161
      8181 ,    // 8162
      8181 ,    // 8163
      8181 ,    // 8164
      8181 ,    // 8165
      8181 ,    // 8166
      8181 ,    // 8167
      8181 ,    // 8168
      8181 ,    // 8169
      8181 ,    // 8170
      8181 ,    // 8171
      8181 ,    // 8172
      8181 ,    // 8173
      8181 ,    // 8174
      8181 ,    // 8175
      8181 ,    // 8176
      8181 ,    // 8177
      8181 ,    // 8178
      8181 ,    // 8179
      8181 ,    // 8180
      8181 ,    // 8181
      8181 ,    // 8182
      8181 ,    // 8183
      8181 ,    // 8184
      8181 ,    // 8185
      8181 ,    // 8186
      8181 ,    // 8187
      8181 ,    // 8188

      8181 ,    // 8189
      8181 ,    // 8190
      8181      // 8191
};

  logic [12:0] iadr0_;
  logic [12:0] iadr1_;

  always_ff @(posedge iclk) begin
    if (iclkena) begin
      iadr0_ <= iadr0;
      odat0  <= coe[iadr0_];

      iadr1_ <= iadr1;
      odat1  <= coe[iadr1_];
    end
  end
endmodule